library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"64440000",
     1 => x"444c5c74",
     2 => x"08080000",
     3 => x"4141773e",
     4 => x"00000000",
     5 => x"00007f7f",
     6 => x"41410000",
     7 => x"08083e77",
     8 => x"01010200",
     9 => x"01020203",
    10 => x"7f7f7f00",
    11 => x"7f7f7f7f",
    12 => x"1c080800",
    13 => x"7f3e3e1c",
    14 => x"3e7f7f7f",
    15 => x"081c1c3e",
    16 => x"18100008",
    17 => x"10187c7c",
    18 => x"30100000",
    19 => x"10307c7c",
    20 => x"60301000",
    21 => x"061e7860",
    22 => x"3c664200",
    23 => x"42663c18",
    24 => x"6a387800",
    25 => x"386cc6c2",
    26 => x"00006000",
    27 => x"60000060",
    28 => x"5b5e0e00",
    29 => x"1e0e5d5c",
    30 => x"eec24c71",
    31 => x"c04dbfdd",
    32 => x"741ec04b",
    33 => x"87c702ab",
    34 => x"c048a6c4",
    35 => x"c487c578",
    36 => x"78c148a6",
    37 => x"731e66c4",
    38 => x"87dfee49",
    39 => x"e0c086c8",
    40 => x"87eeef49",
    41 => x"6a4aa5c4",
    42 => x"87f0f049",
    43 => x"cb87c6f1",
    44 => x"c883c185",
    45 => x"ff04abb7",
    46 => x"262687c7",
    47 => x"264c264d",
    48 => x"1e4f264b",
    49 => x"eec24a71",
    50 => x"eec25ae1",
    51 => x"78c748e1",
    52 => x"87ddfe49",
    53 => x"731e4f26",
    54 => x"c04a711e",
    55 => x"d303aab7",
    56 => x"d8d3c287",
    57 => x"87c405bf",
    58 => x"87c24bc1",
    59 => x"d3c24bc0",
    60 => x"87c45bdc",
    61 => x"5adcd3c2",
    62 => x"bfd8d3c2",
    63 => x"c19ac14a",
    64 => x"ec49a2c0",
    65 => x"48fc87e8",
    66 => x"bfd8d3c2",
    67 => x"87effe78",
    68 => x"c44a711e",
    69 => x"49721e66",
    70 => x"2687f9ea",
    71 => x"ff1e4f26",
    72 => x"ffc348d4",
    73 => x"48d0ff78",
    74 => x"ff78e1c0",
    75 => x"78c148d4",
    76 => x"30c44871",
    77 => x"7808d4ff",
    78 => x"c048d0ff",
    79 => x"4f2678e0",
    80 => x"5c5b5e0e",
    81 => x"86f40e5d",
    82 => x"c048a6c4",
    83 => x"bfec4b78",
    84 => x"ddeec27e",
    85 => x"bfe84dbf",
    86 => x"d8d3c24c",
    87 => x"fee249bf",
    88 => x"49eecb87",
    89 => x"cc87f9cd",
    90 => x"49c758a6",
    91 => x"7087f3e6",
    92 => x"87c80598",
    93 => x"99c1496e",
    94 => x"87c3c102",
    95 => x"bfec4bc1",
    96 => x"d8d3c27e",
    97 => x"d6e249bf",
    98 => x"4966c887",
    99 => x"7087ddcd",
   100 => x"87d80298",
   101 => x"bfc0d3c2",
   102 => x"c2b9c149",
   103 => x"7159c4d3",
   104 => x"cb87fbfd",
   105 => x"f7cc49ee",
   106 => x"58a6cc87",
   107 => x"f1e549c7",
   108 => x"05987087",
   109 => x"6e87c5ff",
   110 => x"0599c149",
   111 => x"7387fdfe",
   112 => x"87d0029b",
   113 => x"cdfc49ff",
   114 => x"49dac187",
   115 => x"c487d3e5",
   116 => x"78c148a6",
   117 => x"bfd8d3c2",
   118 => x"87d9c105",
   119 => x"c848a6c4",
   120 => x"c278c0c0",
   121 => x"6e7ec4d3",
   122 => x"6e49bf97",
   123 => x"7080c148",
   124 => x"ede4717e",
   125 => x"02987087",
   126 => x"66c487c3",
   127 => x"4866c4b4",
   128 => x"c828b7c1",
   129 => x"987058a6",
   130 => x"87dbff05",
   131 => x"e449fdc3",
   132 => x"fac387d0",
   133 => x"87cae449",
   134 => x"ffc34974",
   135 => x"c01e7199",
   136 => x"87ecfb49",
   137 => x"b7c84974",
   138 => x"c11e7129",
   139 => x"87e0fb49",
   140 => x"f4c886c8",
   141 => x"c3497487",
   142 => x"b7c899ff",
   143 => x"74b4712c",
   144 => x"87df029c",
   145 => x"bfd4d3c2",
   146 => x"87e0ca49",
   147 => x"c0059870",
   148 => x"4cc087c4",
   149 => x"e0c287d3",
   150 => x"87c4ca49",
   151 => x"58d8d3c2",
   152 => x"c287c6c0",
   153 => x"c048d4d3",
   154 => x"c2497478",
   155 => x"cec00599",
   156 => x"49ebc387",
   157 => x"7087ebe2",
   158 => x"0299c249",
   159 => x"c187cfc0",
   160 => x"6e7ea5d8",
   161 => x"c5c002bf",
   162 => x"49fb4b87",
   163 => x"49740f73",
   164 => x"c00599c1",
   165 => x"f4c387ce",
   166 => x"87c6e249",
   167 => x"99c24970",
   168 => x"87cfc002",
   169 => x"7ea5d8c1",
   170 => x"c002bf6e",
   171 => x"fa4b87c5",
   172 => x"740f7349",
   173 => x"0599c849",
   174 => x"c387cec0",
   175 => x"e1e149f5",
   176 => x"c2497087",
   177 => x"e5c00299",
   178 => x"e1eec287",
   179 => x"cac002bf",
   180 => x"88c14887",
   181 => x"58e5eec2",
   182 => x"c187cec0",
   183 => x"6a4aa5d8",
   184 => x"87c5c002",
   185 => x"7349ff4b",
   186 => x"48a6c40f",
   187 => x"497478c1",
   188 => x"c00599c4",
   189 => x"f2c387ce",
   190 => x"87e6e049",
   191 => x"99c24970",
   192 => x"87ecc002",
   193 => x"bfe1eec2",
   194 => x"b7c7487e",
   195 => x"cbc003a8",
   196 => x"c1486e87",
   197 => x"e5eec280",
   198 => x"87cfc058",
   199 => x"7ea5d8c1",
   200 => x"c002bf6e",
   201 => x"fe4b87c5",
   202 => x"c40f7349",
   203 => x"78c148a6",
   204 => x"ff49fdc3",
   205 => x"7087ebdf",
   206 => x"0299c249",
   207 => x"c287e5c0",
   208 => x"02bfe1ee",
   209 => x"c287c9c0",
   210 => x"c048e1ee",
   211 => x"87cfc078",
   212 => x"7ea5d8c1",
   213 => x"c002bf6e",
   214 => x"fd4b87c5",
   215 => x"c40f7349",
   216 => x"78c148a6",
   217 => x"ff49fac3",
   218 => x"7087f7de",
   219 => x"0299c249",
   220 => x"c287e9c0",
   221 => x"48bfe1ee",
   222 => x"03a8b7c7",
   223 => x"c287c9c0",
   224 => x"c748e1ee",
   225 => x"87cfc078",
   226 => x"7ea5d8c1",
   227 => x"c002bf6e",
   228 => x"fc4b87c5",
   229 => x"c40f7349",
   230 => x"78c148a6",
   231 => x"eec24bc0",
   232 => x"50c048dc",
   233 => x"c449eecb",
   234 => x"a6cc87f6",
   235 => x"dceec258",
   236 => x"c105bf97",
   237 => x"497487de",
   238 => x"0599f0c3",
   239 => x"c187cdc0",
   240 => x"ddff49da",
   241 => x"987087dc",
   242 => x"87c8c102",
   243 => x"bfe84bc1",
   244 => x"ffc3494c",
   245 => x"2cb7c899",
   246 => x"d3c2b471",
   247 => x"ff49bfd8",
   248 => x"c887fcd8",
   249 => x"c3c44966",
   250 => x"02987087",
   251 => x"c287c6c0",
   252 => x"c148dcee",
   253 => x"dceec250",
   254 => x"c005bf97",
   255 => x"497487d6",
   256 => x"0599f0c3",
   257 => x"c187c5ff",
   258 => x"dcff49da",
   259 => x"987087d4",
   260 => x"87f8fe05",
   261 => x"c0029b73",
   262 => x"a6c887dc",
   263 => x"e1eec248",
   264 => x"66c878bf",
   265 => x"7591cb49",
   266 => x"bf6e7ea1",
   267 => x"87c6c002",
   268 => x"4966c84b",
   269 => x"66c40f73",
   270 => x"87c8c002",
   271 => x"bfe1eec2",
   272 => x"87edf049",
   273 => x"bfdcd3c2",
   274 => x"87ddc002",
   275 => x"87dcc249",
   276 => x"c0029870",
   277 => x"eec287d3",
   278 => x"f049bfe1",
   279 => x"49c087d3",
   280 => x"c287f3f1",
   281 => x"c048dcd3",
   282 => x"f18ef478",
   283 => x"5e0e87cd",
   284 => x"0e5d5c5b",
   285 => x"c24c711e",
   286 => x"49bfddee",
   287 => x"4da1cdc1",
   288 => x"6981d1c1",
   289 => x"029c747e",
   290 => x"a5c487cf",
   291 => x"c27b744b",
   292 => x"49bfddee",
   293 => x"6e87ecf0",
   294 => x"059c747b",
   295 => x"4bc087c4",
   296 => x"4bc187c2",
   297 => x"edf04973",
   298 => x"0266d487",
   299 => x"c04987c8",
   300 => x"4a7087ee",
   301 => x"4ac087c2",
   302 => x"5ae0d3c2",
   303 => x"87fbef26",
   304 => x"00000000",
   305 => x"14111258",
   306 => x"231c1b1d",
   307 => x"9491595a",
   308 => x"f4ebf2f5",
   309 => x"00000000",
   310 => x"00000000",
   311 => x"00000000",
   312 => x"ff4a711e",
   313 => x"7249bfc8",
   314 => x"4f2648a1",
   315 => x"bfc8ff1e",
   316 => x"c0c0fe89",
   317 => x"a9c0c0c0",
   318 => x"c087c401",
   319 => x"c187c24a",
   320 => x"2648724a",
   321 => x"5b5e0e4f",
   322 => x"710e5d5c",
   323 => x"4cd4ff4b",
   324 => x"c04866d0",
   325 => x"ff49d678",
   326 => x"c387ffd9",
   327 => x"496c7cff",
   328 => x"7199ffc3",
   329 => x"f0c3494d",
   330 => x"a9e0c199",
   331 => x"c387cb05",
   332 => x"486c7cff",
   333 => x"66d098c3",
   334 => x"ffc37808",
   335 => x"494a6c7c",
   336 => x"ffc331c8",
   337 => x"714a6c7c",
   338 => x"c84972b2",
   339 => x"7cffc331",
   340 => x"b2714a6c",
   341 => x"31c84972",
   342 => x"6c7cffc3",
   343 => x"ffb2714a",
   344 => x"e0c048d0",
   345 => x"029b7378",
   346 => x"7b7287c2",
   347 => x"4d264875",
   348 => x"4b264c26",
   349 => x"261e4f26",
   350 => x"5b5e0e4f",
   351 => x"86f80e5c",
   352 => x"a6c81e76",
   353 => x"87fdfd49",
   354 => x"4b7086c4",
   355 => x"a8c2486e",
   356 => x"87f0c203",
   357 => x"f0c34a73",
   358 => x"aad0c19a",
   359 => x"c187c702",
   360 => x"c205aae0",
   361 => x"497387de",
   362 => x"c30299c8",
   363 => x"87c6ff87",
   364 => x"9cc34c73",
   365 => x"c105acc2",
   366 => x"66c487c2",
   367 => x"7131c949",
   368 => x"4a66c41e",
   369 => x"eec292d4",
   370 => x"817249e5",
   371 => x"87f7cffe",
   372 => x"d7ff49d8",
   373 => x"c0c887c4",
   374 => x"ceddc21e",
   375 => x"fdebfd49",
   376 => x"48d0ff87",
   377 => x"c278e0c0",
   378 => x"cc1ecedd",
   379 => x"92d44a66",
   380 => x"49e5eec2",
   381 => x"cdfe8172",
   382 => x"86cc87ff",
   383 => x"c105acc1",
   384 => x"66c487c2",
   385 => x"7131c949",
   386 => x"4a66c41e",
   387 => x"eec292d4",
   388 => x"817249e5",
   389 => x"87efcefe",
   390 => x"1eceddc2",
   391 => x"d44a66c8",
   392 => x"e5eec292",
   393 => x"fe817249",
   394 => x"d787c0cc",
   395 => x"e9d5ff49",
   396 => x"1ec0c887",
   397 => x"49ceddc2",
   398 => x"87fbe9fd",
   399 => x"d0ff86cc",
   400 => x"78e0c048",
   401 => x"e7fc8ef8",
   402 => x"5b5e0e87",
   403 => x"710e5d5c",
   404 => x"4cd4ff4a",
   405 => x"c34d66d0",
   406 => x"c506adb7",
   407 => x"c148c087",
   408 => x"1e7287e1",
   409 => x"93d44b75",
   410 => x"83e5eec2",
   411 => x"c6fe4973",
   412 => x"83c887c7",
   413 => x"d0ff4b6b",
   414 => x"78e1c848",
   415 => x"48737cdd",
   416 => x"7098ffc3",
   417 => x"c849737c",
   418 => x"487129b7",
   419 => x"7098ffc3",
   420 => x"d049737c",
   421 => x"487129b7",
   422 => x"7098ffc3",
   423 => x"d848737c",
   424 => x"7c7028b7",
   425 => x"7c7c7cc0",
   426 => x"7c7c7c7c",
   427 => x"7c7c7c7c",
   428 => x"48d0ff7c",
   429 => x"7578e0c0",
   430 => x"ff49dc1e",
   431 => x"c887c0d4",
   432 => x"fa487386",
   433 => x"731e87e8",
   434 => x"1e4bc01e",
   435 => x"bfc7dcc2",
   436 => x"87f5fd49",
   437 => x"dcc286c4",
   438 => x"fe49bfcb",
   439 => x"7087d0dd",
   440 => x"87c40598",
   441 => x"4bf4dbc2",
   442 => x"87c44873",
   443 => x"4c264d26",
   444 => x"4f264b26",
   445 => x"204d4f52",
   446 => x"64616f6c",
   447 => x"20676e69",
   448 => x"6c696166",
   449 => x"0f006465",
   450 => x"1b000027",
   451 => x"42000027",
   452 => x"20204342",
   453 => x"56202020",
   454 => x"42004448",
   455 => x"20204342",
   456 => x"52202020",
   457 => x"52004d4f",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
