library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"ccefc287",
    12 => x"86c0c84e",
    13 => x"49ccefc2",
    14 => x"48d8dcc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087fbe1",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d40299",
    50 => x"d4ff4812",
    51 => x"66c47808",
    52 => x"88c14849",
    53 => x"7158a6c8",
    54 => x"87ec0599",
    55 => x"711e4f26",
    56 => x"4966c44a",
    57 => x"c888c148",
    58 => x"997158a6",
    59 => x"ff87d602",
    60 => x"ffc348d4",
    61 => x"c4526878",
    62 => x"c1484966",
    63 => x"58a6c888",
    64 => x"ea059971",
    65 => x"1e4f2687",
    66 => x"d4ff1e73",
    67 => x"7bffc34b",
    68 => x"ffc34a6b",
    69 => x"c8496b7b",
    70 => x"c3b17232",
    71 => x"4a6b7bff",
    72 => x"b27131c8",
    73 => x"6b7bffc3",
    74 => x"7232c849",
    75 => x"c44871b1",
    76 => x"264d2687",
    77 => x"264b264c",
    78 => x"5b5e0e4f",
    79 => x"710e5d5c",
    80 => x"4cd4ff4a",
    81 => x"ffc34872",
    82 => x"c27c7098",
    83 => x"05bfd8dc",
    84 => x"66d087c8",
    85 => x"d430c948",
    86 => x"66d058a6",
    87 => x"7129d849",
    88 => x"98ffc348",
    89 => x"66d07c70",
    90 => x"7129d049",
    91 => x"98ffc348",
    92 => x"66d07c70",
    93 => x"7129c849",
    94 => x"98ffc348",
    95 => x"66d07c70",
    96 => x"98ffc348",
    97 => x"49727c70",
    98 => x"487129d0",
    99 => x"7098ffc3",
   100 => x"c94b6c7c",
   101 => x"c34dfff0",
   102 => x"d005abff",
   103 => x"7cffc387",
   104 => x"8dc14b6c",
   105 => x"c387c602",
   106 => x"f002abff",
   107 => x"fd487387",
   108 => x"c01e87ff",
   109 => x"48d4ff49",
   110 => x"c178ffc3",
   111 => x"b7c8c381",
   112 => x"87f104a9",
   113 => x"731e4f26",
   114 => x"c487e71e",
   115 => x"c04bdff8",
   116 => x"f0ffc01e",
   117 => x"fd49f7c1",
   118 => x"86c487df",
   119 => x"c005a8c1",
   120 => x"d4ff87ea",
   121 => x"78ffc348",
   122 => x"c0c0c0c1",
   123 => x"c01ec0c0",
   124 => x"e9c1f0e1",
   125 => x"87c1fd49",
   126 => x"987086c4",
   127 => x"ff87ca05",
   128 => x"ffc348d4",
   129 => x"cb48c178",
   130 => x"87e6fe87",
   131 => x"fe058bc1",
   132 => x"48c087fd",
   133 => x"1e87defc",
   134 => x"d4ff1e73",
   135 => x"78ffc348",
   136 => x"1ec04bd3",
   137 => x"c1f0ffc0",
   138 => x"ccfc49c1",
   139 => x"7086c487",
   140 => x"87ca0598",
   141 => x"c348d4ff",
   142 => x"48c178ff",
   143 => x"f1fd87cb",
   144 => x"058bc187",
   145 => x"c087dbff",
   146 => x"87e9fb48",
   147 => x"5c5b5e0e",
   148 => x"4cd4ff0e",
   149 => x"c687dbfd",
   150 => x"e1c01eea",
   151 => x"49c8c1f0",
   152 => x"c487d6fb",
   153 => x"02a8c186",
   154 => x"eafe87c8",
   155 => x"c148c087",
   156 => x"d2fa87e2",
   157 => x"cf497087",
   158 => x"c699ffff",
   159 => x"c802a9ea",
   160 => x"87d3fe87",
   161 => x"cbc148c0",
   162 => x"7cffc387",
   163 => x"fc4bf1c0",
   164 => x"987087f4",
   165 => x"87ebc002",
   166 => x"ffc01ec0",
   167 => x"49fac1f0",
   168 => x"c487d6fa",
   169 => x"05987086",
   170 => x"ffc387d9",
   171 => x"c3496c7c",
   172 => x"7c7c7cff",
   173 => x"99c0c17c",
   174 => x"c187c402",
   175 => x"c087d548",
   176 => x"c287d148",
   177 => x"87c405ab",
   178 => x"87c848c0",
   179 => x"fe058bc1",
   180 => x"48c087fd",
   181 => x"1e87dcf9",
   182 => x"dcc21e73",
   183 => x"78c148d8",
   184 => x"d0ff4bc7",
   185 => x"fb78c248",
   186 => x"d0ff87c8",
   187 => x"c078c348",
   188 => x"d0e5c01e",
   189 => x"f849c0c1",
   190 => x"86c487ff",
   191 => x"c105a8c1",
   192 => x"abc24b87",
   193 => x"c087c505",
   194 => x"87f9c048",
   195 => x"ff058bc1",
   196 => x"f7fc87d0",
   197 => x"dcdcc287",
   198 => x"05987058",
   199 => x"1ec187cd",
   200 => x"c1f0ffc0",
   201 => x"d0f849d0",
   202 => x"ff86c487",
   203 => x"ffc348d4",
   204 => x"87ddc478",
   205 => x"58e0dcc2",
   206 => x"c248d0ff",
   207 => x"48d4ff78",
   208 => x"c178ffc3",
   209 => x"87edf748",
   210 => x"5c5b5e0e",
   211 => x"4a710e5d",
   212 => x"ff4dffc3",
   213 => x"7c754cd4",
   214 => x"c448d0ff",
   215 => x"7c7578c3",
   216 => x"ffc01e72",
   217 => x"49d8c1f0",
   218 => x"c487cef7",
   219 => x"02987086",
   220 => x"48c187c5",
   221 => x"7587eec0",
   222 => x"7cfec37c",
   223 => x"d41ec0c8",
   224 => x"f2f44966",
   225 => x"7586c487",
   226 => x"757c757c",
   227 => x"e0dad87c",
   228 => x"6c7c754b",
   229 => x"c187c505",
   230 => x"87f5058b",
   231 => x"d0ff7c75",
   232 => x"c078c248",
   233 => x"87c9f648",
   234 => x"5c5b5e0e",
   235 => x"4b710e5d",
   236 => x"eec54cc0",
   237 => x"ff4adfcd",
   238 => x"ffc348d4",
   239 => x"c3486878",
   240 => x"c005a8fe",
   241 => x"d4ff87fe",
   242 => x"029b734d",
   243 => x"66d087cc",
   244 => x"f449731e",
   245 => x"86c487c8",
   246 => x"d0ff87d6",
   247 => x"78d1c448",
   248 => x"d07dffc3",
   249 => x"88c14866",
   250 => x"7058a6d4",
   251 => x"87f00598",
   252 => x"c348d4ff",
   253 => x"737878ff",
   254 => x"87c5059b",
   255 => x"d048d0ff",
   256 => x"4c4ac178",
   257 => x"fe058ac1",
   258 => x"487487ed",
   259 => x"1e87e2f4",
   260 => x"4a711e73",
   261 => x"d4ff4bc0",
   262 => x"78ffc348",
   263 => x"c448d0ff",
   264 => x"d4ff78c3",
   265 => x"78ffc348",
   266 => x"ffc01e72",
   267 => x"49d1c1f0",
   268 => x"c487c6f4",
   269 => x"05987086",
   270 => x"c0c887d2",
   271 => x"4966cc1e",
   272 => x"c487e5fd",
   273 => x"ff4b7086",
   274 => x"78c248d0",
   275 => x"e4f34873",
   276 => x"5b5e0e87",
   277 => x"c00e5d5c",
   278 => x"f0ffc01e",
   279 => x"f349c9c1",
   280 => x"1ed287d7",
   281 => x"49e0dcc2",
   282 => x"c887fdfc",
   283 => x"c14cc086",
   284 => x"acb7d284",
   285 => x"c287f804",
   286 => x"bf97e0dc",
   287 => x"99c0c349",
   288 => x"05a9c0c1",
   289 => x"c287e7c0",
   290 => x"bf97e7dc",
   291 => x"c231d049",
   292 => x"bf97e8dc",
   293 => x"7232c84a",
   294 => x"e9dcc2b1",
   295 => x"b14abf97",
   296 => x"ffcf4c71",
   297 => x"c19cffff",
   298 => x"c134ca84",
   299 => x"dcc287e7",
   300 => x"49bf97e9",
   301 => x"99c631c1",
   302 => x"97eadcc2",
   303 => x"b7c74abf",
   304 => x"c2b1722a",
   305 => x"bf97e5dc",
   306 => x"9dcf4d4a",
   307 => x"97e6dcc2",
   308 => x"9ac34abf",
   309 => x"dcc232ca",
   310 => x"4bbf97e7",
   311 => x"b27333c2",
   312 => x"97e8dcc2",
   313 => x"c0c34bbf",
   314 => x"2bb7c69b",
   315 => x"81c2b273",
   316 => x"307148c1",
   317 => x"48c14970",
   318 => x"4d703075",
   319 => x"84c14c72",
   320 => x"c0c89471",
   321 => x"cc06adb7",
   322 => x"b734c187",
   323 => x"b7c0c82d",
   324 => x"f4ff01ad",
   325 => x"f0487487",
   326 => x"5e0e87d7",
   327 => x"0e5d5c5b",
   328 => x"e5c286f8",
   329 => x"78c048c6",
   330 => x"1efedcc2",
   331 => x"defb49c0",
   332 => x"7086c487",
   333 => x"87c50598",
   334 => x"c0c948c0",
   335 => x"c14dc087",
   336 => x"ddf2c07e",
   337 => x"ddc249bf",
   338 => x"c8714af4",
   339 => x"87d9ec4b",
   340 => x"c2059870",
   341 => x"c07ec087",
   342 => x"49bfd9f2",
   343 => x"4ad0dec2",
   344 => x"ec4bc871",
   345 => x"987087c3",
   346 => x"c087c205",
   347 => x"c0026e7e",
   348 => x"e4c287fd",
   349 => x"c24dbfc4",
   350 => x"bf9ffce4",
   351 => x"d6c5487e",
   352 => x"c705a8ea",
   353 => x"c4e4c287",
   354 => x"87ce4dbf",
   355 => x"e9ca486e",
   356 => x"c502a8d5",
   357 => x"c748c087",
   358 => x"dcc287e3",
   359 => x"49751efe",
   360 => x"c487ecf9",
   361 => x"05987086",
   362 => x"48c087c5",
   363 => x"c087cec7",
   364 => x"49bfd9f2",
   365 => x"4ad0dec2",
   366 => x"ea4bc871",
   367 => x"987087eb",
   368 => x"c287c805",
   369 => x"c148c6e5",
   370 => x"c087da78",
   371 => x"49bfddf2",
   372 => x"4af4ddc2",
   373 => x"ea4bc871",
   374 => x"987087cf",
   375 => x"87c5c002",
   376 => x"d8c648c0",
   377 => x"fce4c287",
   378 => x"c149bf97",
   379 => x"c005a9d5",
   380 => x"e4c287cd",
   381 => x"49bf97fd",
   382 => x"02a9eac2",
   383 => x"c087c5c0",
   384 => x"87f9c548",
   385 => x"97fedcc2",
   386 => x"c3487ebf",
   387 => x"c002a8e9",
   388 => x"486e87ce",
   389 => x"02a8ebc3",
   390 => x"c087c5c0",
   391 => x"87ddc548",
   392 => x"97c9ddc2",
   393 => x"059949bf",
   394 => x"c287ccc0",
   395 => x"bf97cadd",
   396 => x"02a9c249",
   397 => x"c087c5c0",
   398 => x"87c1c548",
   399 => x"97cbddc2",
   400 => x"e5c248bf",
   401 => x"4c7058c2",
   402 => x"c288c148",
   403 => x"c258c6e5",
   404 => x"bf97ccdd",
   405 => x"c2817549",
   406 => x"bf97cddd",
   407 => x"7232c84a",
   408 => x"e9c27ea1",
   409 => x"786e48d3",
   410 => x"97ceddc2",
   411 => x"a6c848bf",
   412 => x"c6e5c258",
   413 => x"cfc202bf",
   414 => x"d9f2c087",
   415 => x"dec249bf",
   416 => x"c8714ad0",
   417 => x"87e1e74b",
   418 => x"c0029870",
   419 => x"48c087c5",
   420 => x"c287eac3",
   421 => x"4cbffee4",
   422 => x"5ce7e9c2",
   423 => x"97e3ddc2",
   424 => x"31c849bf",
   425 => x"97e2ddc2",
   426 => x"49a14abf",
   427 => x"97e4ddc2",
   428 => x"32d04abf",
   429 => x"c249a172",
   430 => x"bf97e5dd",
   431 => x"7232d84a",
   432 => x"66c449a1",
   433 => x"d3e9c291",
   434 => x"e9c281bf",
   435 => x"ddc259db",
   436 => x"4abf97eb",
   437 => x"ddc232c8",
   438 => x"4bbf97ea",
   439 => x"ddc24aa2",
   440 => x"4bbf97ec",
   441 => x"a27333d0",
   442 => x"edddc24a",
   443 => x"cf4bbf97",
   444 => x"7333d89b",
   445 => x"e9c24aa2",
   446 => x"8ac25adf",
   447 => x"e9c29274",
   448 => x"a17248df",
   449 => x"87c1c178",
   450 => x"97d0ddc2",
   451 => x"31c849bf",
   452 => x"97cfddc2",
   453 => x"49a14abf",
   454 => x"ffc731c5",
   455 => x"c229c981",
   456 => x"c259e7e9",
   457 => x"bf97d5dd",
   458 => x"c232c84a",
   459 => x"bf97d4dd",
   460 => x"c44aa24b",
   461 => x"826e9266",
   462 => x"5ae3e9c2",
   463 => x"48dbe9c2",
   464 => x"e9c278c0",
   465 => x"a17248d7",
   466 => x"e7e9c278",
   467 => x"dbe9c248",
   468 => x"e9c278bf",
   469 => x"e9c248eb",
   470 => x"c278bfdf",
   471 => x"02bfc6e5",
   472 => x"7487c9c0",
   473 => x"7030c448",
   474 => x"87c9c07e",
   475 => x"bfe3e9c2",
   476 => x"7030c448",
   477 => x"cae5c27e",
   478 => x"c1786e48",
   479 => x"268ef848",
   480 => x"264c264d",
   481 => x"0e4f264b",
   482 => x"5d5c5b5e",
   483 => x"c24a710e",
   484 => x"02bfc6e5",
   485 => x"4b7287cb",
   486 => x"4d722bc7",
   487 => x"c99dffc1",
   488 => x"c84b7287",
   489 => x"c34d722b",
   490 => x"e9c29dff",
   491 => x"c083bfd3",
   492 => x"abbfd5f2",
   493 => x"c087d902",
   494 => x"c25bd9f2",
   495 => x"731efedc",
   496 => x"87cbf149",
   497 => x"987086c4",
   498 => x"c087c505",
   499 => x"87e6c048",
   500 => x"bfc6e5c2",
   501 => x"7587d202",
   502 => x"c291c449",
   503 => x"6981fedc",
   504 => x"ffffcf4c",
   505 => x"cb9cffff",
   506 => x"c2497587",
   507 => x"fedcc291",
   508 => x"4c699f81",
   509 => x"c6fe4874",
   510 => x"5b5e0e87",
   511 => x"f80e5d5c",
   512 => x"9c4c7186",
   513 => x"c087c505",
   514 => x"87c0c348",
   515 => x"487ea4c8",
   516 => x"66d878c0",
   517 => x"d887c702",
   518 => x"05bf9766",
   519 => x"48c087c5",
   520 => x"c087e9c2",
   521 => x"4949c11e",
   522 => x"c487d3ca",
   523 => x"9d4d7086",
   524 => x"87c2c102",
   525 => x"4acee5c2",
   526 => x"e04966d8",
   527 => x"987087d0",
   528 => x"87f2c002",
   529 => x"66d84a75",
   530 => x"e04bcb49",
   531 => x"987087f5",
   532 => x"87e2c002",
   533 => x"9d751ec0",
   534 => x"c887c702",
   535 => x"78c048a6",
   536 => x"a6c887c5",
   537 => x"c878c148",
   538 => x"d1c94966",
   539 => x"7086c487",
   540 => x"fe059d4d",
   541 => x"9d7587fe",
   542 => x"87cec102",
   543 => x"6e49a5dc",
   544 => x"da786948",
   545 => x"a6c449a5",
   546 => x"78a4c448",
   547 => x"c448699f",
   548 => x"c2780866",
   549 => x"02bfc6e5",
   550 => x"a5d487d2",
   551 => x"49699f49",
   552 => x"99ffffc0",
   553 => x"30d04871",
   554 => x"87c27e70",
   555 => x"486e7ec0",
   556 => x"80bf66c4",
   557 => x"780866c4",
   558 => x"a4cc7cc0",
   559 => x"bf66c449",
   560 => x"49a4d079",
   561 => x"48c179c0",
   562 => x"48c087c2",
   563 => x"eefa8ef8",
   564 => x"5b5e0e87",
   565 => x"4c710e5c",
   566 => x"cbc1029c",
   567 => x"49a4c887",
   568 => x"c3c10269",
   569 => x"cc496c87",
   570 => x"80714866",
   571 => x"7058a6d0",
   572 => x"c2e5c2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e5c002",
   576 => x"6b4ba4c4",
   577 => x"87fff949",
   578 => x"e4c27b70",
   579 => x"6c49bffe",
   580 => x"cc7c7181",
   581 => x"e5c2b966",
   582 => x"ff4abfc2",
   583 => x"719972ba",
   584 => x"dbff0599",
   585 => x"7c66cc87",
   586 => x"1e87d6f9",
   587 => x"4b711e73",
   588 => x"87c7029b",
   589 => x"6949a3c8",
   590 => x"c087c505",
   591 => x"87f6c048",
   592 => x"bfd7e9c2",
   593 => x"4aa3c449",
   594 => x"8ac24a6a",
   595 => x"bffee4c2",
   596 => x"49a17292",
   597 => x"bfc2e5c2",
   598 => x"729a6b4a",
   599 => x"f2c049a1",
   600 => x"66c859d9",
   601 => x"e6ea711e",
   602 => x"7086c487",
   603 => x"87c40598",
   604 => x"87c248c0",
   605 => x"caf848c1",
   606 => x"1e731e87",
   607 => x"029b4b71",
   608 => x"a3c887c7",
   609 => x"c5056949",
   610 => x"c048c087",
   611 => x"e9c287f6",
   612 => x"c449bfd7",
   613 => x"4a6a4aa3",
   614 => x"e4c28ac2",
   615 => x"7292bffe",
   616 => x"e5c249a1",
   617 => x"6b4abfc2",
   618 => x"49a1729a",
   619 => x"59d9f2c0",
   620 => x"711e66c8",
   621 => x"c487d1e6",
   622 => x"05987086",
   623 => x"48c087c4",
   624 => x"48c187c2",
   625 => x"0e87fcf6",
   626 => x"5d5c5b5e",
   627 => x"4b711e0e",
   628 => x"734d66d4",
   629 => x"ccc1029b",
   630 => x"49a3c887",
   631 => x"c4c10269",
   632 => x"4ca3d087",
   633 => x"bfc2e5c2",
   634 => x"6cb9ff49",
   635 => x"d47e994a",
   636 => x"cd06a966",
   637 => x"7c7bc087",
   638 => x"c44aa3cc",
   639 => x"796a49a3",
   640 => x"497287ca",
   641 => x"d499c0f8",
   642 => x"8d714d66",
   643 => x"29c94975",
   644 => x"49731e71",
   645 => x"c287fafa",
   646 => x"731efedc",
   647 => x"87cbfc49",
   648 => x"66d486c8",
   649 => x"d6f5267c",
   650 => x"1e731e87",
   651 => x"029b4b71",
   652 => x"c287e4c0",
   653 => x"735bebe9",
   654 => x"c28ac24a",
   655 => x"49bffee4",
   656 => x"d7e9c292",
   657 => x"807248bf",
   658 => x"58efe9c2",
   659 => x"30c44871",
   660 => x"58cee5c2",
   661 => x"c287edc0",
   662 => x"c248e7e9",
   663 => x"78bfdbe9",
   664 => x"48ebe9c2",
   665 => x"bfdfe9c2",
   666 => x"c6e5c278",
   667 => x"87c902bf",
   668 => x"bffee4c2",
   669 => x"c731c449",
   670 => x"e3e9c287",
   671 => x"31c449bf",
   672 => x"59cee5c2",
   673 => x"0e87fcf3",
   674 => x"0e5c5b5e",
   675 => x"4bc04a71",
   676 => x"c0029a72",
   677 => x"a2da87e0",
   678 => x"4b699f49",
   679 => x"bfc6e5c2",
   680 => x"d487cf02",
   681 => x"699f49a2",
   682 => x"ffc04c49",
   683 => x"34d09cff",
   684 => x"4cc087c2",
   685 => x"4973b374",
   686 => x"f387eefd",
   687 => x"5e0e87c3",
   688 => x"0e5d5c5b",
   689 => x"4a7186f4",
   690 => x"9a727ec0",
   691 => x"c287d802",
   692 => x"c048fadc",
   693 => x"f2dcc278",
   694 => x"ebe9c248",
   695 => x"dcc278bf",
   696 => x"e9c248f6",
   697 => x"c278bfe7",
   698 => x"c048dbe5",
   699 => x"cae5c250",
   700 => x"dcc249bf",
   701 => x"714abffa",
   702 => x"c9c403aa",
   703 => x"cf497287",
   704 => x"e9c00599",
   705 => x"d5f2c087",
   706 => x"f2dcc248",
   707 => x"dcc278bf",
   708 => x"dcc21efe",
   709 => x"c249bff2",
   710 => x"c148f2dc",
   711 => x"e37178a1",
   712 => x"86c487ed",
   713 => x"48d1f2c0",
   714 => x"78fedcc2",
   715 => x"f2c087cc",
   716 => x"c048bfd1",
   717 => x"f2c080e0",
   718 => x"dcc258d5",
   719 => x"c148bffa",
   720 => x"fedcc280",
   721 => x"0c912758",
   722 => x"97bf0000",
   723 => x"029d4dbf",
   724 => x"c387e3c2",
   725 => x"c202ade5",
   726 => x"f2c087dc",
   727 => x"cb4bbfd1",
   728 => x"4c1149a3",
   729 => x"c105accf",
   730 => x"497587d2",
   731 => x"89c199df",
   732 => x"e5c291cd",
   733 => x"a3c181ce",
   734 => x"c351124a",
   735 => x"51124aa3",
   736 => x"124aa3c5",
   737 => x"4aa3c751",
   738 => x"a3c95112",
   739 => x"ce51124a",
   740 => x"51124aa3",
   741 => x"124aa3d0",
   742 => x"4aa3d251",
   743 => x"a3d45112",
   744 => x"d651124a",
   745 => x"51124aa3",
   746 => x"124aa3d8",
   747 => x"4aa3dc51",
   748 => x"a3de5112",
   749 => x"c151124a",
   750 => x"87fac07e",
   751 => x"99c84974",
   752 => x"87ebc005",
   753 => x"99d04974",
   754 => x"dc87d105",
   755 => x"cbc00266",
   756 => x"dc497387",
   757 => x"98700f66",
   758 => x"87d3c002",
   759 => x"c6c0056e",
   760 => x"cee5c287",
   761 => x"c050c048",
   762 => x"48bfd1f2",
   763 => x"c287ddc2",
   764 => x"c048dbe5",
   765 => x"e5c27e50",
   766 => x"c249bfca",
   767 => x"4abffadc",
   768 => x"fb04aa71",
   769 => x"e9c287f7",
   770 => x"c005bfeb",
   771 => x"e5c287c8",
   772 => x"c102bfc6",
   773 => x"dcc287f4",
   774 => x"ed49bff6",
   775 => x"dcc287e9",
   776 => x"a6c458fa",
   777 => x"f6dcc248",
   778 => x"e5c278bf",
   779 => x"c002bfc6",
   780 => x"66c487d8",
   781 => x"ffffcf49",
   782 => x"a999f8ff",
   783 => x"87c5c002",
   784 => x"e1c04cc0",
   785 => x"c04cc187",
   786 => x"66c487dc",
   787 => x"f8ffcf49",
   788 => x"c002a999",
   789 => x"a6c887c8",
   790 => x"c078c048",
   791 => x"a6c887c5",
   792 => x"c878c148",
   793 => x"9c744c66",
   794 => x"87dec005",
   795 => x"c24966c4",
   796 => x"fee4c289",
   797 => x"e9c291bf",
   798 => x"7148bfd7",
   799 => x"f6dcc280",
   800 => x"fadcc258",
   801 => x"f978c048",
   802 => x"48c087e3",
   803 => x"eeeb8ef4",
   804 => x"00000087",
   805 => x"ffffff00",
   806 => x"000ca1ff",
   807 => x"000caa00",
   808 => x"54414600",
   809 => x"20203233",
   810 => x"41460020",
   811 => x"20363154",
   812 => x"1e002020",
   813 => x"c348d4ff",
   814 => x"486878ff",
   815 => x"ff1e4f26",
   816 => x"ffc348d4",
   817 => x"48d0ff78",
   818 => x"ff78e1c0",
   819 => x"78d448d4",
   820 => x"48efe9c2",
   821 => x"50bfd4ff",
   822 => x"ff1e4f26",
   823 => x"e0c048d0",
   824 => x"1e4f2678",
   825 => x"7087ccff",
   826 => x"c6029949",
   827 => x"a9fbc087",
   828 => x"7187f105",
   829 => x"0e4f2648",
   830 => x"0e5c5b5e",
   831 => x"4cc04b71",
   832 => x"7087f0fe",
   833 => x"c0029949",
   834 => x"ecc087f9",
   835 => x"f2c002a9",
   836 => x"a9fbc087",
   837 => x"87ebc002",
   838 => x"acb766cc",
   839 => x"d087c703",
   840 => x"87c20266",
   841 => x"99715371",
   842 => x"c187c202",
   843 => x"87c3fe84",
   844 => x"02994970",
   845 => x"ecc087cd",
   846 => x"87c702a9",
   847 => x"05a9fbc0",
   848 => x"d087d5ff",
   849 => x"87c30266",
   850 => x"c07b97c0",
   851 => x"c405a9ec",
   852 => x"c54a7487",
   853 => x"c04a7487",
   854 => x"48728a0a",
   855 => x"4d2687c2",
   856 => x"4b264c26",
   857 => x"fd1e4f26",
   858 => x"497087c9",
   859 => x"aaf0c04a",
   860 => x"c087c904",
   861 => x"c301aaf9",
   862 => x"8af0c087",
   863 => x"04aac1c1",
   864 => x"dac187c9",
   865 => x"87c301aa",
   866 => x"728af7c0",
   867 => x"0e4f2648",
   868 => x"0e5c5b5e",
   869 => x"d4ff4a71",
   870 => x"c049724b",
   871 => x"4c7087e7",
   872 => x"87c2029c",
   873 => x"d0ff8cc1",
   874 => x"c178c548",
   875 => x"49747bd5",
   876 => x"e3c131c6",
   877 => x"4abf97dc",
   878 => x"70b07148",
   879 => x"48d0ff7b",
   880 => x"dbfe78c4",
   881 => x"5b5e0e87",
   882 => x"f80e5d5c",
   883 => x"c04c7186",
   884 => x"87eafb7e",
   885 => x"f9c04bc0",
   886 => x"49bf97f2",
   887 => x"cf04a9c0",
   888 => x"87fffb87",
   889 => x"f9c083c1",
   890 => x"49bf97f2",
   891 => x"87f106ab",
   892 => x"97f2f9c0",
   893 => x"87cf02bf",
   894 => x"7087f8fa",
   895 => x"c6029949",
   896 => x"a9ecc087",
   897 => x"c087f105",
   898 => x"87e7fa4b",
   899 => x"e2fa4d70",
   900 => x"58a6c887",
   901 => x"7087dcfa",
   902 => x"c883c14a",
   903 => x"699749a4",
   904 => x"c702ad49",
   905 => x"adffc087",
   906 => x"87e7c005",
   907 => x"9749a4c9",
   908 => x"66c44969",
   909 => x"87c702a9",
   910 => x"a8ffc048",
   911 => x"ca87d405",
   912 => x"699749a4",
   913 => x"c602aa49",
   914 => x"aaffc087",
   915 => x"c187c405",
   916 => x"c087d07e",
   917 => x"c602adec",
   918 => x"adfbc087",
   919 => x"c087c405",
   920 => x"6e7ec14b",
   921 => x"87e1fe02",
   922 => x"7387eff9",
   923 => x"fb8ef848",
   924 => x"0e0087ec",
   925 => x"5d5c5b5e",
   926 => x"7186f80e",
   927 => x"4bd4ff4d",
   928 => x"e9c21e75",
   929 => x"f0e549f4",
   930 => x"7086c487",
   931 => x"cac40298",
   932 => x"48a6c487",
   933 => x"bfdee3c1",
   934 => x"fb497578",
   935 => x"d0ff87f1",
   936 => x"c178c548",
   937 => x"4ac07bd6",
   938 => x"1149a275",
   939 => x"cb82c17b",
   940 => x"f304aab7",
   941 => x"c34acc87",
   942 => x"82c17bff",
   943 => x"aab7e0c0",
   944 => x"ff87f404",
   945 => x"78c448d0",
   946 => x"c57bffc3",
   947 => x"7bd3c178",
   948 => x"78c47bc1",
   949 => x"b7c04866",
   950 => x"eec206a8",
   951 => x"fce9c287",
   952 => x"66c44cbf",
   953 => x"c8887448",
   954 => x"9c7458a6",
   955 => x"87f7c102",
   956 => x"7efedcc2",
   957 => x"8c4dc0c8",
   958 => x"03acb7c0",
   959 => x"c0c887c6",
   960 => x"4cc04da4",
   961 => x"97efe9c2",
   962 => x"99d049bf",
   963 => x"c087d002",
   964 => x"f4e9c21e",
   965 => x"87d3e849",
   966 => x"4a7086c4",
   967 => x"c287edc0",
   968 => x"c21efedc",
   969 => x"e849f4e9",
   970 => x"86c487c1",
   971 => x"d0ff4a70",
   972 => x"78c5c848",
   973 => x"6e7bd4c1",
   974 => x"6e7bbf97",
   975 => x"7080c148",
   976 => x"058dc17e",
   977 => x"ff87f0ff",
   978 => x"78c448d0",
   979 => x"c5059a72",
   980 => x"c148c087",
   981 => x"1ec187c7",
   982 => x"49f4e9c2",
   983 => x"c487f2e5",
   984 => x"059c7486",
   985 => x"c487c9fe",
   986 => x"b7c04866",
   987 => x"87d106a8",
   988 => x"48f4e9c2",
   989 => x"80d078c0",
   990 => x"80f478c0",
   991 => x"bfc0eac2",
   992 => x"4866c478",
   993 => x"01a8b7c0",
   994 => x"ff87d2fd",
   995 => x"78c548d0",
   996 => x"c07bd3c1",
   997 => x"c178c47b",
   998 => x"c087c248",
   999 => x"268ef848",
  1000 => x"264c264d",
  1001 => x"0e4f264b",
  1002 => x"5d5c5b5e",
  1003 => x"4b711e0e",
  1004 => x"ab4d4cc0",
  1005 => x"87e8c004",
  1006 => x"1ec5f7c0",
  1007 => x"c4029d75",
  1008 => x"c24ac087",
  1009 => x"724ac187",
  1010 => x"87f2eb49",
  1011 => x"7e7086c4",
  1012 => x"056e84c1",
  1013 => x"4c7387c2",
  1014 => x"ac7385c1",
  1015 => x"87d8ff06",
  1016 => x"fe26486e",
  1017 => x"5e0e87f9",
  1018 => x"710e5c5b",
  1019 => x"0266cc4b",
  1020 => x"c04c87d8",
  1021 => x"d8028cf0",
  1022 => x"c14a7487",
  1023 => x"87d1028a",
  1024 => x"87cd028a",
  1025 => x"87c9028a",
  1026 => x"497387d9",
  1027 => x"d287e4f9",
  1028 => x"c01e7487",
  1029 => x"d6d8c149",
  1030 => x"731e7487",
  1031 => x"ced8c149",
  1032 => x"fd86c887",
  1033 => x"5e0e87fb",
  1034 => x"0e5d5c5b",
  1035 => x"494c711e",
  1036 => x"eac291de",
  1037 => x"85714ddc",
  1038 => x"c1026d97",
  1039 => x"eac287dc",
  1040 => x"7449bfc8",
  1041 => x"defd7181",
  1042 => x"487e7087",
  1043 => x"f2c00298",
  1044 => x"d0eac287",
  1045 => x"cb4a704b",
  1046 => x"cac1ff49",
  1047 => x"cb4b7487",
  1048 => x"f0e3c193",
  1049 => x"c183c483",
  1050 => x"747bdec2",
  1051 => x"e5c0c149",
  1052 => x"c17b7587",
  1053 => x"bf97dde3",
  1054 => x"eac21e49",
  1055 => x"e5fd49d0",
  1056 => x"7486c487",
  1057 => x"cdc0c149",
  1058 => x"c149c087",
  1059 => x"c287ecc1",
  1060 => x"c048f0e9",
  1061 => x"dd49c178",
  1062 => x"fc2687fb",
  1063 => x"6f4c87c1",
  1064 => x"6e696461",
  1065 => x"2e2e2e67",
  1066 => x"1e731e00",
  1067 => x"c2494a71",
  1068 => x"81bfc8ea",
  1069 => x"87effb71",
  1070 => x"029b4b70",
  1071 => x"e74987c4",
  1072 => x"eac287c5",
  1073 => x"78c048c8",
  1074 => x"c8dd49c1",
  1075 => x"87d3fb87",
  1076 => x"5c5b5e0e",
  1077 => x"86f40e5d",
  1078 => x"4dfedcc2",
  1079 => x"a6c44cc0",
  1080 => x"c278c048",
  1081 => x"48bfc8ea",
  1082 => x"c106a8c0",
  1083 => x"dcc287c0",
  1084 => x"029848fe",
  1085 => x"c087f7c0",
  1086 => x"c81ec5f7",
  1087 => x"87c70266",
  1088 => x"c048a6c4",
  1089 => x"c487c578",
  1090 => x"78c148a6",
  1091 => x"e64966c4",
  1092 => x"86c487ec",
  1093 => x"84c14d70",
  1094 => x"c14866c4",
  1095 => x"58a6c880",
  1096 => x"bfc8eac2",
  1097 => x"87c603ac",
  1098 => x"ff059d75",
  1099 => x"4cc087c9",
  1100 => x"c3029d75",
  1101 => x"f7c087dc",
  1102 => x"66c81ec5",
  1103 => x"cc87c702",
  1104 => x"78c048a6",
  1105 => x"a6cc87c5",
  1106 => x"cc78c148",
  1107 => x"ede54966",
  1108 => x"7086c487",
  1109 => x"0298487e",
  1110 => x"4987e4c2",
  1111 => x"699781cb",
  1112 => x"0299d049",
  1113 => x"7487d4c1",
  1114 => x"c191cb49",
  1115 => x"c181f0e3",
  1116 => x"c879e9c2",
  1117 => x"51ffc381",
  1118 => x"91de4974",
  1119 => x"4ddceac2",
  1120 => x"c1c28571",
  1121 => x"a5c17d97",
  1122 => x"51e0c049",
  1123 => x"97cee5c2",
  1124 => x"87d202bf",
  1125 => x"a5c284c1",
  1126 => x"cee5c24b",
  1127 => x"fe49db4a",
  1128 => x"c187c4fc",
  1129 => x"a5cd87d9",
  1130 => x"c151c049",
  1131 => x"4ba5c284",
  1132 => x"49cb4a6e",
  1133 => x"87effbfe",
  1134 => x"7487c4c1",
  1135 => x"c191cb49",
  1136 => x"c181f0e3",
  1137 => x"c279e6c0",
  1138 => x"bf97cee5",
  1139 => x"7487d802",
  1140 => x"c191de49",
  1141 => x"dceac284",
  1142 => x"c283714b",
  1143 => x"dd4acee5",
  1144 => x"c2fbfe49",
  1145 => x"7487d887",
  1146 => x"c293de4b",
  1147 => x"cb83dcea",
  1148 => x"51c049a3",
  1149 => x"6e7384c1",
  1150 => x"fe49cb4a",
  1151 => x"c487e8fa",
  1152 => x"80c14866",
  1153 => x"c758a6c8",
  1154 => x"c5c003ac",
  1155 => x"fc056e87",
  1156 => x"487487e4",
  1157 => x"c6f68ef4",
  1158 => x"1e731e87",
  1159 => x"cb494b71",
  1160 => x"f0e3c191",
  1161 => x"4aa1c881",
  1162 => x"48dce3c1",
  1163 => x"a1c95012",
  1164 => x"f2f9c04a",
  1165 => x"ca501248",
  1166 => x"dde3c181",
  1167 => x"c1501148",
  1168 => x"bf97dde3",
  1169 => x"49c01e49",
  1170 => x"c287dbf6",
  1171 => x"de48f0e9",
  1172 => x"d649c178",
  1173 => x"f52687ff",
  1174 => x"711e87c9",
  1175 => x"91cb494a",
  1176 => x"81f0e3c1",
  1177 => x"481181c8",
  1178 => x"58f4e9c2",
  1179 => x"48c8eac2",
  1180 => x"49c178c0",
  1181 => x"2687ded6",
  1182 => x"49c01e4f",
  1183 => x"87fbf9c0",
  1184 => x"711e4f26",
  1185 => x"87d20299",
  1186 => x"48c5e5c1",
  1187 => x"80f750c0",
  1188 => x"40dac9c1",
  1189 => x"78e9e3c1",
  1190 => x"e5c187ce",
  1191 => x"e3c148c1",
  1192 => x"80fc78e2",
  1193 => x"78f9c9c1",
  1194 => x"5e0e4f26",
  1195 => x"0e5d5c5b",
  1196 => x"4d7186f4",
  1197 => x"c191cb49",
  1198 => x"c881f0e3",
  1199 => x"a1ca4aa1",
  1200 => x"48a6c47e",
  1201 => x"bff8edc2",
  1202 => x"bf976e78",
  1203 => x"4c66c44b",
  1204 => x"48122c73",
  1205 => x"7058a6cc",
  1206 => x"c984c19c",
  1207 => x"49699781",
  1208 => x"c204acb7",
  1209 => x"6e4cc087",
  1210 => x"c84abf97",
  1211 => x"31724966",
  1212 => x"66c4b9ff",
  1213 => x"72487499",
  1214 => x"484a7030",
  1215 => x"edc2b071",
  1216 => x"e4c058fc",
  1217 => x"49c087d0",
  1218 => x"7587cad4",
  1219 => x"c5f6c049",
  1220 => x"f28ef487",
  1221 => x"731e87c9",
  1222 => x"494b711e",
  1223 => x"7387cbfe",
  1224 => x"87c6fe49",
  1225 => x"1e87fcf1",
  1226 => x"4b711e73",
  1227 => x"024aa3c6",
  1228 => x"8ac187db",
  1229 => x"8a87d602",
  1230 => x"87dac102",
  1231 => x"fcc0028a",
  1232 => x"c0028a87",
  1233 => x"028a87e1",
  1234 => x"dbc187cb",
  1235 => x"fc49c787",
  1236 => x"dec187c8",
  1237 => x"c8eac287",
  1238 => x"cbc102bf",
  1239 => x"88c14887",
  1240 => x"58cceac2",
  1241 => x"c287c1c1",
  1242 => x"02bfccea",
  1243 => x"c287f9c0",
  1244 => x"48bfc8ea",
  1245 => x"eac280c1",
  1246 => x"ebc058cc",
  1247 => x"c8eac287",
  1248 => x"89c649bf",
  1249 => x"59cceac2",
  1250 => x"03a9b7c0",
  1251 => x"eac287da",
  1252 => x"78c048c8",
  1253 => x"eac287d2",
  1254 => x"cb02bfcc",
  1255 => x"c8eac287",
  1256 => x"80c648bf",
  1257 => x"58cceac2",
  1258 => x"e8d149c0",
  1259 => x"c0497387",
  1260 => x"ef87e3f3",
  1261 => x"5e0e87ed",
  1262 => x"0e5d5c5b",
  1263 => x"dc86d4ff",
  1264 => x"a6c859a6",
  1265 => x"c478c048",
  1266 => x"66c0c180",
  1267 => x"c180c478",
  1268 => x"c180c478",
  1269 => x"cceac278",
  1270 => x"c278c148",
  1271 => x"48bff0e9",
  1272 => x"c905a8de",
  1273 => x"87e8f387",
  1274 => x"cf58a6cc",
  1275 => x"cde387e6",
  1276 => x"87efe387",
  1277 => x"7087fce2",
  1278 => x"acfbc04c",
  1279 => x"87fbc102",
  1280 => x"c10566d8",
  1281 => x"fcc087ed",
  1282 => x"82c44a66",
  1283 => x"1e727e6a",
  1284 => x"48c9e0c1",
  1285 => x"c84966c4",
  1286 => x"41204aa1",
  1287 => x"f905aa71",
  1288 => x"26511087",
  1289 => x"66fcc04a",
  1290 => x"d9c8c148",
  1291 => x"c7496a78",
  1292 => x"c0517481",
  1293 => x"c84966fc",
  1294 => x"c051c181",
  1295 => x"c94966fc",
  1296 => x"c051c081",
  1297 => x"ca4966fc",
  1298 => x"c151c081",
  1299 => x"6a1ed81e",
  1300 => x"e281c849",
  1301 => x"86c887e1",
  1302 => x"4866c0c1",
  1303 => x"c701a8c0",
  1304 => x"48a6c887",
  1305 => x"87ce78c1",
  1306 => x"4866c0c1",
  1307 => x"a6d088c1",
  1308 => x"e187c358",
  1309 => x"a6d087ed",
  1310 => x"7478c248",
  1311 => x"cfcd029c",
  1312 => x"4866c887",
  1313 => x"a866c4c1",
  1314 => x"87c4cd03",
  1315 => x"c048a6dc",
  1316 => x"c080e878",
  1317 => x"87dbe078",
  1318 => x"d0c14c70",
  1319 => x"d7c205ac",
  1320 => x"7e66c487",
  1321 => x"c887ffe2",
  1322 => x"c6e058a6",
  1323 => x"c04c7087",
  1324 => x"c105acec",
  1325 => x"66c887ed",
  1326 => x"c091cb49",
  1327 => x"c48166fc",
  1328 => x"4d6a4aa1",
  1329 => x"c44aa1c8",
  1330 => x"c9c15266",
  1331 => x"dfff79da",
  1332 => x"4c7087e1",
  1333 => x"87d9029c",
  1334 => x"02acfbc0",
  1335 => x"557487d3",
  1336 => x"87cfdfff",
  1337 => x"029c4c70",
  1338 => x"fbc087c7",
  1339 => x"edff05ac",
  1340 => x"55e0c087",
  1341 => x"c055c1c2",
  1342 => x"66d87d97",
  1343 => x"05a86e48",
  1344 => x"66c887db",
  1345 => x"a866cc48",
  1346 => x"c887ca04",
  1347 => x"80c14866",
  1348 => x"c858a6cc",
  1349 => x"4866cc87",
  1350 => x"a6d088c1",
  1351 => x"d2deff58",
  1352 => x"c14c7087",
  1353 => x"c805acd0",
  1354 => x"4866d487",
  1355 => x"a6d880c1",
  1356 => x"acd0c158",
  1357 => x"87e9fd02",
  1358 => x"d84866c4",
  1359 => x"c905a866",
  1360 => x"e0c087e0",
  1361 => x"78c048a6",
  1362 => x"fbc04874",
  1363 => x"487e7088",
  1364 => x"e2c90298",
  1365 => x"88cb4887",
  1366 => x"98487e70",
  1367 => x"87cdc102",
  1368 => x"7088c948",
  1369 => x"0298487e",
  1370 => x"4887fec3",
  1371 => x"7e7088c4",
  1372 => x"ce029848",
  1373 => x"88c14887",
  1374 => x"98487e70",
  1375 => x"87e9c302",
  1376 => x"dc87d6c8",
  1377 => x"f0c048a6",
  1378 => x"e6dcff78",
  1379 => x"c04c7087",
  1380 => x"c002acec",
  1381 => x"e0c087c4",
  1382 => x"ecc05ca6",
  1383 => x"87cd02ac",
  1384 => x"87cfdcff",
  1385 => x"ecc04c70",
  1386 => x"f3ff05ac",
  1387 => x"acecc087",
  1388 => x"87c4c002",
  1389 => x"87fbdbff",
  1390 => x"1eca1ec0",
  1391 => x"cb4966d0",
  1392 => x"66c4c191",
  1393 => x"cc807148",
  1394 => x"66c858a6",
  1395 => x"d080c448",
  1396 => x"66cc58a6",
  1397 => x"dcff49bf",
  1398 => x"1ec187dd",
  1399 => x"66d41ede",
  1400 => x"dcff49bf",
  1401 => x"86d087d1",
  1402 => x"c0484970",
  1403 => x"e8c08808",
  1404 => x"a8c058a6",
  1405 => x"87eec006",
  1406 => x"4866e4c0",
  1407 => x"c003a8dd",
  1408 => x"66c487e4",
  1409 => x"e4c049bf",
  1410 => x"e0c08166",
  1411 => x"66e4c051",
  1412 => x"c481c149",
  1413 => x"c281bf66",
  1414 => x"e4c051c1",
  1415 => x"81c24966",
  1416 => x"81bf66c4",
  1417 => x"486e51c0",
  1418 => x"78d9c8c1",
  1419 => x"81c8496e",
  1420 => x"6e5166d0",
  1421 => x"d481c949",
  1422 => x"496e5166",
  1423 => x"66dc81ca",
  1424 => x"4866d051",
  1425 => x"a6d480c1",
  1426 => x"4866c858",
  1427 => x"04a866cc",
  1428 => x"c887cbc0",
  1429 => x"80c14866",
  1430 => x"c558a6cc",
  1431 => x"66cc87d9",
  1432 => x"d088c148",
  1433 => x"cec558a6",
  1434 => x"f9dbff87",
  1435 => x"a6e8c087",
  1436 => x"f1dbff58",
  1437 => x"a6e0c087",
  1438 => x"a8ecc058",
  1439 => x"87cac005",
  1440 => x"c048a6dc",
  1441 => x"c07866e4",
  1442 => x"d8ff87c4",
  1443 => x"66c887e5",
  1444 => x"c091cb49",
  1445 => x"714866fc",
  1446 => x"4a7e7080",
  1447 => x"496e82c8",
  1448 => x"e4c081ca",
  1449 => x"66dc5166",
  1450 => x"c081c149",
  1451 => x"c18966e4",
  1452 => x"70307148",
  1453 => x"7189c149",
  1454 => x"edc27a97",
  1455 => x"c049bff8",
  1456 => x"972966e4",
  1457 => x"71484a6a",
  1458 => x"a6ecc098",
  1459 => x"c4496e58",
  1460 => x"d84d6981",
  1461 => x"66c44866",
  1462 => x"c8c002a8",
  1463 => x"48a6c487",
  1464 => x"c5c078c0",
  1465 => x"48a6c487",
  1466 => x"66c478c1",
  1467 => x"1ee0c01e",
  1468 => x"d8ff4975",
  1469 => x"86c887c1",
  1470 => x"b7c04c70",
  1471 => x"d4c106ac",
  1472 => x"c0857487",
  1473 => x"897449e0",
  1474 => x"e0c14b75",
  1475 => x"fe714ad2",
  1476 => x"c287d4e6",
  1477 => x"66e0c085",
  1478 => x"c080c148",
  1479 => x"c058a6e4",
  1480 => x"c14966e8",
  1481 => x"02a97081",
  1482 => x"c487c8c0",
  1483 => x"78c048a6",
  1484 => x"c487c5c0",
  1485 => x"78c148a6",
  1486 => x"c21e66c4",
  1487 => x"e0c049a4",
  1488 => x"70887148",
  1489 => x"49751e49",
  1490 => x"87ebd6ff",
  1491 => x"b7c086c8",
  1492 => x"c0ff01a8",
  1493 => x"66e0c087",
  1494 => x"87d1c002",
  1495 => x"81c9496e",
  1496 => x"5166e0c0",
  1497 => x"cac1486e",
  1498 => x"ccc078ea",
  1499 => x"c9496e87",
  1500 => x"6e51c281",
  1501 => x"d6ccc148",
  1502 => x"4866c878",
  1503 => x"04a866cc",
  1504 => x"c887cbc0",
  1505 => x"80c14866",
  1506 => x"c058a6cc",
  1507 => x"66cc87e9",
  1508 => x"d088c148",
  1509 => x"dec058a6",
  1510 => x"c6d5ff87",
  1511 => x"c04c7087",
  1512 => x"c6c187d5",
  1513 => x"c8c005ac",
  1514 => x"4866d087",
  1515 => x"a6d480c1",
  1516 => x"eed4ff58",
  1517 => x"d44c7087",
  1518 => x"80c14866",
  1519 => x"7458a6d8",
  1520 => x"cbc0029c",
  1521 => x"4866c887",
  1522 => x"a866c4c1",
  1523 => x"87fcf204",
  1524 => x"87c6d4ff",
  1525 => x"c74866c8",
  1526 => x"e5c003a8",
  1527 => x"cceac287",
  1528 => x"c878c048",
  1529 => x"91cb4966",
  1530 => x"8166fcc0",
  1531 => x"6a4aa1c4",
  1532 => x"7952c04a",
  1533 => x"c14866c8",
  1534 => x"58a6cc80",
  1535 => x"ff04a8c7",
  1536 => x"d4ff87db",
  1537 => x"d6deff8e",
  1538 => x"616f4c87",
  1539 => x"2e2a2064",
  1540 => x"203a0020",
  1541 => x"1e731e00",
  1542 => x"029b4b71",
  1543 => x"eac287c6",
  1544 => x"78c048c8",
  1545 => x"eac21ec7",
  1546 => x"c11ebfc8",
  1547 => x"c21ef0e3",
  1548 => x"49bff0e9",
  1549 => x"cc87ffed",
  1550 => x"f0e9c286",
  1551 => x"c1e949bf",
  1552 => x"029b7387",
  1553 => x"e3c187c8",
  1554 => x"e2c049f0",
  1555 => x"ddff87da",
  1556 => x"c71e87d1",
  1557 => x"49c187d1",
  1558 => x"fe87fafe",
  1559 => x"7087f8e9",
  1560 => x"87cd0298",
  1561 => x"87f2f2fe",
  1562 => x"c4029870",
  1563 => x"c24ac187",
  1564 => x"724ac087",
  1565 => x"87ce059a",
  1566 => x"e2c11ec0",
  1567 => x"efc049e3",
  1568 => x"86c487d2",
  1569 => x"1ec087fe",
  1570 => x"49eee2c1",
  1571 => x"87c4efc0",
  1572 => x"f8c01ec0",
  1573 => x"497087e1",
  1574 => x"87f8eec0",
  1575 => x"f887c7c3",
  1576 => x"534f268e",
  1577 => x"61662044",
  1578 => x"64656c69",
  1579 => x"6f42002e",
  1580 => x"6e69746f",
  1581 => x"2e2e2e67",
  1582 => x"e5c01e00",
  1583 => x"f2c087e7",
  1584 => x"87f687dd",
  1585 => x"c21e4f26",
  1586 => x"c048c8ea",
  1587 => x"f0e9c278",
  1588 => x"fd78c048",
  1589 => x"87e187fc",
  1590 => x"4f2648c0",
  1591 => x"00010000",
  1592 => x"20800000",
  1593 => x"74697845",
  1594 => x"42208000",
  1595 => x"006b6361",
  1596 => x"00001026",
  1597 => x"00002a9c",
  1598 => x"26000000",
  1599 => x"ba000010",
  1600 => x"0000002a",
  1601 => x"10260000",
  1602 => x"2ad80000",
  1603 => x"00000000",
  1604 => x"00102600",
  1605 => x"002af600",
  1606 => x"00000000",
  1607 => x"00001026",
  1608 => x"00002b14",
  1609 => x"26000000",
  1610 => x"32000010",
  1611 => x"0000002b",
  1612 => x"10260000",
  1613 => x"2b500000",
  1614 => x"00000000",
  1615 => x"00125a00",
  1616 => x"00000000",
  1617 => x"00000000",
  1618 => x"00001327",
  1619 => x"00000000",
  1620 => x"1e000000",
  1621 => x"c048f0fe",
  1622 => x"7909cd78",
  1623 => x"1e4f2609",
  1624 => x"48bff0fe",
  1625 => x"fe1e4f26",
  1626 => x"78c148f0",
  1627 => x"fe1e4f26",
  1628 => x"78c048f0",
  1629 => x"711e4f26",
  1630 => x"5152c04a",
  1631 => x"5e0e4f26",
  1632 => x"0e5d5c5b",
  1633 => x"4d7186f4",
  1634 => x"c17e6d97",
  1635 => x"6c974ca5",
  1636 => x"58a6c848",
  1637 => x"66c4486e",
  1638 => x"87c505a8",
  1639 => x"e6c048ff",
  1640 => x"87caff87",
  1641 => x"9749a5c2",
  1642 => x"a3714b6c",
  1643 => x"4b6b974b",
  1644 => x"6e7e6c97",
  1645 => x"c880c148",
  1646 => x"98c758a6",
  1647 => x"7058a6cc",
  1648 => x"e1fe7c97",
  1649 => x"f4487387",
  1650 => x"264d268e",
  1651 => x"264b264c",
  1652 => x"5b5e0e4f",
  1653 => x"86f40e5c",
  1654 => x"66d84c71",
  1655 => x"9affc34a",
  1656 => x"974ba4c2",
  1657 => x"a173496c",
  1658 => x"97517249",
  1659 => x"486e7e6c",
  1660 => x"a6c880c1",
  1661 => x"cc98c758",
  1662 => x"547058a6",
  1663 => x"caff8ef4",
  1664 => x"fd1e1e87",
  1665 => x"bfe087e8",
  1666 => x"e0c0494a",
  1667 => x"cb0299c0",
  1668 => x"c21e7287",
  1669 => x"fe49eeed",
  1670 => x"86c487f7",
  1671 => x"7087c0fd",
  1672 => x"87c2fd7e",
  1673 => x"1e4f2626",
  1674 => x"49eeedc2",
  1675 => x"c187c7fd",
  1676 => x"fc49c1e8",
  1677 => x"f7c387dd",
  1678 => x"0e4f2687",
  1679 => x"5d5c5b5e",
  1680 => x"c24d710e",
  1681 => x"fc49eeed",
  1682 => x"4b7087f4",
  1683 => x"04abb7c0",
  1684 => x"c387c2c3",
  1685 => x"c905abf0",
  1686 => x"dfecc187",
  1687 => x"c278c148",
  1688 => x"e0c387e3",
  1689 => x"87c905ab",
  1690 => x"48e3ecc1",
  1691 => x"d4c278c1",
  1692 => x"e3ecc187",
  1693 => x"87c602bf",
  1694 => x"4ca3c0c2",
  1695 => x"4c7387c2",
  1696 => x"bfdfecc1",
  1697 => x"87e0c002",
  1698 => x"b7c44974",
  1699 => x"edc19129",
  1700 => x"4a7481ff",
  1701 => x"92c29acf",
  1702 => x"307248c1",
  1703 => x"baff4a70",
  1704 => x"98694872",
  1705 => x"87db7970",
  1706 => x"b7c44974",
  1707 => x"edc19129",
  1708 => x"4a7481ff",
  1709 => x"92c29acf",
  1710 => x"307248c3",
  1711 => x"69484a70",
  1712 => x"757970b0",
  1713 => x"f0c0059d",
  1714 => x"48d0ff87",
  1715 => x"ff78e1c8",
  1716 => x"78c548d4",
  1717 => x"bfe3ecc1",
  1718 => x"c387c302",
  1719 => x"ecc178e0",
  1720 => x"c602bfdf",
  1721 => x"48d4ff87",
  1722 => x"ff78f0c3",
  1723 => x"0b7b0bd4",
  1724 => x"c848d0ff",
  1725 => x"e0c078e1",
  1726 => x"e3ecc178",
  1727 => x"c178c048",
  1728 => x"c048dfec",
  1729 => x"eeedc278",
  1730 => x"87f2f949",
  1731 => x"b7c04b70",
  1732 => x"fefc03ab",
  1733 => x"2648c087",
  1734 => x"264c264d",
  1735 => x"004f264b",
  1736 => x"00000000",
  1737 => x"1e000000",
  1738 => x"fc494a71",
  1739 => x"4f2687cd",
  1740 => x"724ac01e",
  1741 => x"c191c449",
  1742 => x"c081ffed",
  1743 => x"d082c179",
  1744 => x"ee04aab7",
  1745 => x"0e4f2687",
  1746 => x"5d5c5b5e",
  1747 => x"f84d710e",
  1748 => x"4a7587dc",
  1749 => x"922ab7c4",
  1750 => x"82ffedc1",
  1751 => x"9ccf4c75",
  1752 => x"496a94c2",
  1753 => x"c32b744b",
  1754 => x"7448c29b",
  1755 => x"ff4c7030",
  1756 => x"714874bc",
  1757 => x"f77a7098",
  1758 => x"487387ec",
  1759 => x"0087d8fe",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"1e000000",
  1776 => x"c848d0ff",
  1777 => x"487178e1",
  1778 => x"7808d4ff",
  1779 => x"ff1e4f26",
  1780 => x"e1c848d0",
  1781 => x"ff487178",
  1782 => x"c47808d4",
  1783 => x"d4ff4866",
  1784 => x"4f267808",
  1785 => x"c44a711e",
  1786 => x"721e4966",
  1787 => x"87deff49",
  1788 => x"c048d0ff",
  1789 => x"262678e0",
  1790 => x"1e731e4f",
  1791 => x"66c84b71",
  1792 => x"4a731e49",
  1793 => x"49a2e0c1",
  1794 => x"2687d9ff",
  1795 => x"4d2687c4",
  1796 => x"4b264c26",
  1797 => x"ff1e4f26",
  1798 => x"ffc34ad4",
  1799 => x"48d0ff7a",
  1800 => x"de78e1c0",
  1801 => x"f8edc27a",
  1802 => x"48497abf",
  1803 => x"7a7028c8",
  1804 => x"28d04871",
  1805 => x"48717a70",
  1806 => x"7a7028d8",
  1807 => x"c048d0ff",
  1808 => x"4f2678e0",
  1809 => x"48d0ff1e",
  1810 => x"7178c9c8",
  1811 => x"08d4ff48",
  1812 => x"1e4f2678",
  1813 => x"eb494a71",
  1814 => x"48d0ff87",
  1815 => x"4f2678c8",
  1816 => x"711e731e",
  1817 => x"c8eec24b",
  1818 => x"87c302bf",
  1819 => x"ff87ebc2",
  1820 => x"c9c848d0",
  1821 => x"c0487378",
  1822 => x"d4ffb0e0",
  1823 => x"edc27808",
  1824 => x"78c048fc",
  1825 => x"c50266c8",
  1826 => x"49ffc387",
  1827 => x"49c087c2",
  1828 => x"59c4eec2",
  1829 => x"c60266cc",
  1830 => x"d5d5c587",
  1831 => x"cf87c44a",
  1832 => x"c24affff",
  1833 => x"c25ac8ee",
  1834 => x"c148c8ee",
  1835 => x"2687c478",
  1836 => x"264c264d",
  1837 => x"0e4f264b",
  1838 => x"5d5c5b5e",
  1839 => x"c24a710e",
  1840 => x"4cbfc4ee",
  1841 => x"cb029a72",
  1842 => x"91c84987",
  1843 => x"4bd6f1c1",
  1844 => x"87c48371",
  1845 => x"4bd6f5c1",
  1846 => x"49134dc0",
  1847 => x"eec29974",
  1848 => x"7148bfc0",
  1849 => x"08d4ffb8",
  1850 => x"2cb7c178",
  1851 => x"adb7c885",
  1852 => x"c287e704",
  1853 => x"48bffced",
  1854 => x"eec280c8",
  1855 => x"eefe58c0",
  1856 => x"1e731e87",
  1857 => x"4a134b71",
  1858 => x"87cb029a",
  1859 => x"e6fe4972",
  1860 => x"9a4a1387",
  1861 => x"fe87f505",
  1862 => x"c21e87d9",
  1863 => x"49bffced",
  1864 => x"48fcedc2",
  1865 => x"c478a1c1",
  1866 => x"03a9b7c0",
  1867 => x"d4ff87db",
  1868 => x"c0eec248",
  1869 => x"edc278bf",
  1870 => x"c249bffc",
  1871 => x"c148fced",
  1872 => x"c0c478a1",
  1873 => x"e504a9b7",
  1874 => x"48d0ff87",
  1875 => x"eec278c8",
  1876 => x"78c048c8",
  1877 => x"00004f26",
  1878 => x"00000000",
  1879 => x"00000000",
  1880 => x"005f5f00",
  1881 => x"03000000",
  1882 => x"03030003",
  1883 => x"7f140000",
  1884 => x"7f7f147f",
  1885 => x"24000014",
  1886 => x"3a6b6b2e",
  1887 => x"6a4c0012",
  1888 => x"566c1836",
  1889 => x"7e300032",
  1890 => x"3a77594f",
  1891 => x"00004068",
  1892 => x"00030704",
  1893 => x"00000000",
  1894 => x"41633e1c",
  1895 => x"00000000",
  1896 => x"1c3e6341",
  1897 => x"2a080000",
  1898 => x"3e1c1c3e",
  1899 => x"0800082a",
  1900 => x"083e3e08",
  1901 => x"00000008",
  1902 => x"0060e080",
  1903 => x"08000000",
  1904 => x"08080808",
  1905 => x"00000008",
  1906 => x"00606000",
  1907 => x"60400000",
  1908 => x"060c1830",
  1909 => x"3e000103",
  1910 => x"7f4d597f",
  1911 => x"0400003e",
  1912 => x"007f7f06",
  1913 => x"42000000",
  1914 => x"4f597163",
  1915 => x"22000046",
  1916 => x"7f494963",
  1917 => x"1c180036",
  1918 => x"7f7f1316",
  1919 => x"27000010",
  1920 => x"7d454567",
  1921 => x"3c000039",
  1922 => x"79494b7e",
  1923 => x"01000030",
  1924 => x"0f797101",
  1925 => x"36000007",
  1926 => x"7f49497f",
  1927 => x"06000036",
  1928 => x"3f69494f",
  1929 => x"0000001e",
  1930 => x"00666600",
  1931 => x"00000000",
  1932 => x"0066e680",
  1933 => x"08000000",
  1934 => x"22141408",
  1935 => x"14000022",
  1936 => x"14141414",
  1937 => x"22000014",
  1938 => x"08141422",
  1939 => x"02000008",
  1940 => x"0f595103",
  1941 => x"7f3e0006",
  1942 => x"1f555d41",
  1943 => x"7e00001e",
  1944 => x"7f09097f",
  1945 => x"7f00007e",
  1946 => x"7f49497f",
  1947 => x"1c000036",
  1948 => x"4141633e",
  1949 => x"7f000041",
  1950 => x"3e63417f",
  1951 => x"7f00001c",
  1952 => x"4149497f",
  1953 => x"7f000041",
  1954 => x"0109097f",
  1955 => x"3e000001",
  1956 => x"7b49417f",
  1957 => x"7f00007a",
  1958 => x"7f08087f",
  1959 => x"0000007f",
  1960 => x"417f7f41",
  1961 => x"20000000",
  1962 => x"7f404060",
  1963 => x"7f7f003f",
  1964 => x"63361c08",
  1965 => x"7f000041",
  1966 => x"4040407f",
  1967 => x"7f7f0040",
  1968 => x"7f060c06",
  1969 => x"7f7f007f",
  1970 => x"7f180c06",
  1971 => x"3e00007f",
  1972 => x"7f41417f",
  1973 => x"7f00003e",
  1974 => x"0f09097f",
  1975 => x"7f3e0006",
  1976 => x"7e7f6141",
  1977 => x"7f000040",
  1978 => x"7f19097f",
  1979 => x"26000066",
  1980 => x"7b594d6f",
  1981 => x"01000032",
  1982 => x"017f7f01",
  1983 => x"3f000001",
  1984 => x"7f40407f",
  1985 => x"0f00003f",
  1986 => x"3f70703f",
  1987 => x"7f7f000f",
  1988 => x"7f301830",
  1989 => x"6341007f",
  1990 => x"361c1c36",
  1991 => x"03014163",
  1992 => x"067c7c06",
  1993 => x"71610103",
  1994 => x"43474d59",
  1995 => x"00000041",
  1996 => x"41417f7f",
  1997 => x"03010000",
  1998 => x"30180c06",
  1999 => x"00004060",
  2000 => x"7f7f4141",
  2001 => x"0c080000",
  2002 => x"0c060306",
  2003 => x"80800008",
  2004 => x"80808080",
  2005 => x"00000080",
  2006 => x"04070300",
  2007 => x"20000000",
  2008 => x"7c545474",
  2009 => x"7f000078",
  2010 => x"7c44447f",
  2011 => x"38000038",
  2012 => x"4444447c",
  2013 => x"38000000",
  2014 => x"7f44447c",
  2015 => x"3800007f",
  2016 => x"5c54547c",
  2017 => x"04000018",
  2018 => x"05057f7e",
  2019 => x"18000000",
  2020 => x"fca4a4bc",
  2021 => x"7f00007c",
  2022 => x"7c04047f",
  2023 => x"00000078",
  2024 => x"407d3d00",
  2025 => x"80000000",
  2026 => x"7dfd8080",
  2027 => x"7f000000",
  2028 => x"6c38107f",
  2029 => x"00000044",
  2030 => x"407f3f00",
  2031 => x"7c7c0000",
  2032 => x"7c0c180c",
  2033 => x"7c000078",
  2034 => x"7c04047c",
  2035 => x"38000078",
  2036 => x"7c44447c",
  2037 => x"fc000038",
  2038 => x"3c2424fc",
  2039 => x"18000018",
  2040 => x"fc24243c",
  2041 => x"7c0000fc",
  2042 => x"0c04047c",
  2043 => x"48000008",
  2044 => x"7454545c",
  2045 => x"04000020",
  2046 => x"44447f3f",
  2047 => x"3c000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
