
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"cc",x"ef",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"cc",x"ef",x"c2"),
    14 => (x"48",x"d8",x"dc",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"fb",x"e1"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"48",x"72"),
    82 => (x"c2",x"7c",x"70",x"98"),
    83 => (x"05",x"bf",x"d8",x"dc"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"71",x"29",x"d8",x"49"),
    88 => (x"98",x"ff",x"c3",x"48"),
    89 => (x"66",x"d0",x"7c",x"70"),
    90 => (x"71",x"29",x"d0",x"49"),
    91 => (x"98",x"ff",x"c3",x"48"),
    92 => (x"66",x"d0",x"7c",x"70"),
    93 => (x"71",x"29",x"c8",x"49"),
    94 => (x"98",x"ff",x"c3",x"48"),
    95 => (x"66",x"d0",x"7c",x"70"),
    96 => (x"98",x"ff",x"c3",x"48"),
    97 => (x"49",x"72",x"7c",x"70"),
    98 => (x"48",x"71",x"29",x"d0"),
    99 => (x"70",x"98",x"ff",x"c3"),
   100 => (x"c9",x"4b",x"6c",x"7c"),
   101 => (x"c3",x"4d",x"ff",x"f0"),
   102 => (x"d0",x"05",x"ab",x"ff"),
   103 => (x"7c",x"ff",x"c3",x"87"),
   104 => (x"8d",x"c1",x"4b",x"6c"),
   105 => (x"c3",x"87",x"c6",x"02"),
   106 => (x"f0",x"02",x"ab",x"ff"),
   107 => (x"fd",x"48",x"73",x"87"),
   108 => (x"c0",x"1e",x"87",x"ff"),
   109 => (x"48",x"d4",x"ff",x"49"),
   110 => (x"c1",x"78",x"ff",x"c3"),
   111 => (x"b7",x"c8",x"c3",x"81"),
   112 => (x"87",x"f1",x"04",x"a9"),
   113 => (x"73",x"1e",x"4f",x"26"),
   114 => (x"c4",x"87",x"e7",x"1e"),
   115 => (x"c0",x"4b",x"df",x"f8"),
   116 => (x"f0",x"ff",x"c0",x"1e"),
   117 => (x"fd",x"49",x"f7",x"c1"),
   118 => (x"86",x"c4",x"87",x"df"),
   119 => (x"c0",x"05",x"a8",x"c1"),
   120 => (x"d4",x"ff",x"87",x"ea"),
   121 => (x"78",x"ff",x"c3",x"48"),
   122 => (x"c0",x"c0",x"c0",x"c1"),
   123 => (x"c0",x"1e",x"c0",x"c0"),
   124 => (x"e9",x"c1",x"f0",x"e1"),
   125 => (x"87",x"c1",x"fd",x"49"),
   126 => (x"98",x"70",x"86",x"c4"),
   127 => (x"ff",x"87",x"ca",x"05"),
   128 => (x"ff",x"c3",x"48",x"d4"),
   129 => (x"cb",x"48",x"c1",x"78"),
   130 => (x"87",x"e6",x"fe",x"87"),
   131 => (x"fe",x"05",x"8b",x"c1"),
   132 => (x"48",x"c0",x"87",x"fd"),
   133 => (x"1e",x"87",x"de",x"fc"),
   134 => (x"d4",x"ff",x"1e",x"73"),
   135 => (x"78",x"ff",x"c3",x"48"),
   136 => (x"1e",x"c0",x"4b",x"d3"),
   137 => (x"c1",x"f0",x"ff",x"c0"),
   138 => (x"cc",x"fc",x"49",x"c1"),
   139 => (x"70",x"86",x"c4",x"87"),
   140 => (x"87",x"ca",x"05",x"98"),
   141 => (x"c3",x"48",x"d4",x"ff"),
   142 => (x"48",x"c1",x"78",x"ff"),
   143 => (x"f1",x"fd",x"87",x"cb"),
   144 => (x"05",x"8b",x"c1",x"87"),
   145 => (x"c0",x"87",x"db",x"ff"),
   146 => (x"87",x"e9",x"fb",x"48"),
   147 => (x"5c",x"5b",x"5e",x"0e"),
   148 => (x"4c",x"d4",x"ff",x"0e"),
   149 => (x"c6",x"87",x"db",x"fd"),
   150 => (x"e1",x"c0",x"1e",x"ea"),
   151 => (x"49",x"c8",x"c1",x"f0"),
   152 => (x"c4",x"87",x"d6",x"fb"),
   153 => (x"02",x"a8",x"c1",x"86"),
   154 => (x"ea",x"fe",x"87",x"c8"),
   155 => (x"c1",x"48",x"c0",x"87"),
   156 => (x"d2",x"fa",x"87",x"e2"),
   157 => (x"cf",x"49",x"70",x"87"),
   158 => (x"c6",x"99",x"ff",x"ff"),
   159 => (x"c8",x"02",x"a9",x"ea"),
   160 => (x"87",x"d3",x"fe",x"87"),
   161 => (x"cb",x"c1",x"48",x"c0"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"fc",x"4b",x"f1",x"c0"),
   164 => (x"98",x"70",x"87",x"f4"),
   165 => (x"87",x"eb",x"c0",x"02"),
   166 => (x"ff",x"c0",x"1e",x"c0"),
   167 => (x"49",x"fa",x"c1",x"f0"),
   168 => (x"c4",x"87",x"d6",x"fa"),
   169 => (x"05",x"98",x"70",x"86"),
   170 => (x"ff",x"c3",x"87",x"d9"),
   171 => (x"c3",x"49",x"6c",x"7c"),
   172 => (x"7c",x"7c",x"7c",x"ff"),
   173 => (x"99",x"c0",x"c1",x"7c"),
   174 => (x"c1",x"87",x"c4",x"02"),
   175 => (x"c0",x"87",x"d5",x"48"),
   176 => (x"c2",x"87",x"d1",x"48"),
   177 => (x"87",x"c4",x"05",x"ab"),
   178 => (x"87",x"c8",x"48",x"c0"),
   179 => (x"fe",x"05",x"8b",x"c1"),
   180 => (x"48",x"c0",x"87",x"fd"),
   181 => (x"1e",x"87",x"dc",x"f9"),
   182 => (x"dc",x"c2",x"1e",x"73"),
   183 => (x"78",x"c1",x"48",x"d8"),
   184 => (x"d0",x"ff",x"4b",x"c7"),
   185 => (x"fb",x"78",x"c2",x"48"),
   186 => (x"d0",x"ff",x"87",x"c8"),
   187 => (x"c0",x"78",x"c3",x"48"),
   188 => (x"d0",x"e5",x"c0",x"1e"),
   189 => (x"f8",x"49",x"c0",x"c1"),
   190 => (x"86",x"c4",x"87",x"ff"),
   191 => (x"c1",x"05",x"a8",x"c1"),
   192 => (x"ab",x"c2",x"4b",x"87"),
   193 => (x"c0",x"87",x"c5",x"05"),
   194 => (x"87",x"f9",x"c0",x"48"),
   195 => (x"ff",x"05",x"8b",x"c1"),
   196 => (x"f7",x"fc",x"87",x"d0"),
   197 => (x"dc",x"dc",x"c2",x"87"),
   198 => (x"05",x"98",x"70",x"58"),
   199 => (x"1e",x"c1",x"87",x"cd"),
   200 => (x"c1",x"f0",x"ff",x"c0"),
   201 => (x"d0",x"f8",x"49",x"d0"),
   202 => (x"ff",x"86",x"c4",x"87"),
   203 => (x"ff",x"c3",x"48",x"d4"),
   204 => (x"87",x"dd",x"c4",x"78"),
   205 => (x"58",x"e0",x"dc",x"c2"),
   206 => (x"c2",x"48",x"d0",x"ff"),
   207 => (x"48",x"d4",x"ff",x"78"),
   208 => (x"c1",x"78",x"ff",x"c3"),
   209 => (x"87",x"ed",x"f7",x"48"),
   210 => (x"5c",x"5b",x"5e",x"0e"),
   211 => (x"4a",x"71",x"0e",x"5d"),
   212 => (x"ff",x"4d",x"ff",x"c3"),
   213 => (x"7c",x"75",x"4c",x"d4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"7c",x"75",x"78",x"c3"),
   216 => (x"ff",x"c0",x"1e",x"72"),
   217 => (x"49",x"d8",x"c1",x"f0"),
   218 => (x"c4",x"87",x"ce",x"f7"),
   219 => (x"02",x"98",x"70",x"86"),
   220 => (x"48",x"c1",x"87",x"c5"),
   221 => (x"75",x"87",x"ee",x"c0"),
   222 => (x"7c",x"fe",x"c3",x"7c"),
   223 => (x"d4",x"1e",x"c0",x"c8"),
   224 => (x"f2",x"f4",x"49",x"66"),
   225 => (x"75",x"86",x"c4",x"87"),
   226 => (x"75",x"7c",x"75",x"7c"),
   227 => (x"e0",x"da",x"d8",x"7c"),
   228 => (x"6c",x"7c",x"75",x"4b"),
   229 => (x"c1",x"87",x"c5",x"05"),
   230 => (x"87",x"f5",x"05",x"8b"),
   231 => (x"d0",x"ff",x"7c",x"75"),
   232 => (x"c0",x"78",x"c2",x"48"),
   233 => (x"87",x"c9",x"f6",x"48"),
   234 => (x"5c",x"5b",x"5e",x"0e"),
   235 => (x"4b",x"71",x"0e",x"5d"),
   236 => (x"ee",x"c5",x"4c",x"c0"),
   237 => (x"ff",x"4a",x"df",x"cd"),
   238 => (x"ff",x"c3",x"48",x"d4"),
   239 => (x"c3",x"48",x"68",x"78"),
   240 => (x"c0",x"05",x"a8",x"fe"),
   241 => (x"d4",x"ff",x"87",x"fe"),
   242 => (x"02",x"9b",x"73",x"4d"),
   243 => (x"66",x"d0",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c8"),
   246 => (x"d0",x"ff",x"87",x"d6"),
   247 => (x"78",x"d1",x"c4",x"48"),
   248 => (x"d0",x"7d",x"ff",x"c3"),
   249 => (x"88",x"c1",x"48",x"66"),
   250 => (x"70",x"58",x"a6",x"d4"),
   251 => (x"87",x"f0",x"05",x"98"),
   252 => (x"c3",x"48",x"d4",x"ff"),
   253 => (x"73",x"78",x"78",x"ff"),
   254 => (x"87",x"c5",x"05",x"9b"),
   255 => (x"d0",x"48",x"d0",x"ff"),
   256 => (x"4c",x"4a",x"c1",x"78"),
   257 => (x"fe",x"05",x"8a",x"c1"),
   258 => (x"48",x"74",x"87",x"ed"),
   259 => (x"1e",x"87",x"e2",x"f4"),
   260 => (x"4a",x"71",x"1e",x"73"),
   261 => (x"d4",x"ff",x"4b",x"c0"),
   262 => (x"78",x"ff",x"c3",x"48"),
   263 => (x"c4",x"48",x"d0",x"ff"),
   264 => (x"d4",x"ff",x"78",x"c3"),
   265 => (x"78",x"ff",x"c3",x"48"),
   266 => (x"ff",x"c0",x"1e",x"72"),
   267 => (x"49",x"d1",x"c1",x"f0"),
   268 => (x"c4",x"87",x"c6",x"f4"),
   269 => (x"05",x"98",x"70",x"86"),
   270 => (x"c0",x"c8",x"87",x"d2"),
   271 => (x"49",x"66",x"cc",x"1e"),
   272 => (x"c4",x"87",x"e5",x"fd"),
   273 => (x"ff",x"4b",x"70",x"86"),
   274 => (x"78",x"c2",x"48",x"d0"),
   275 => (x"e4",x"f3",x"48",x"73"),
   276 => (x"5b",x"5e",x"0e",x"87"),
   277 => (x"c0",x"0e",x"5d",x"5c"),
   278 => (x"f0",x"ff",x"c0",x"1e"),
   279 => (x"f3",x"49",x"c9",x"c1"),
   280 => (x"1e",x"d2",x"87",x"d7"),
   281 => (x"49",x"e0",x"dc",x"c2"),
   282 => (x"c8",x"87",x"fd",x"fc"),
   283 => (x"c1",x"4c",x"c0",x"86"),
   284 => (x"ac",x"b7",x"d2",x"84"),
   285 => (x"c2",x"87",x"f8",x"04"),
   286 => (x"bf",x"97",x"e0",x"dc"),
   287 => (x"99",x"c0",x"c3",x"49"),
   288 => (x"05",x"a9",x"c0",x"c1"),
   289 => (x"c2",x"87",x"e7",x"c0"),
   290 => (x"bf",x"97",x"e7",x"dc"),
   291 => (x"c2",x"31",x"d0",x"49"),
   292 => (x"bf",x"97",x"e8",x"dc"),
   293 => (x"72",x"32",x"c8",x"4a"),
   294 => (x"e9",x"dc",x"c2",x"b1"),
   295 => (x"b1",x"4a",x"bf",x"97"),
   296 => (x"ff",x"cf",x"4c",x"71"),
   297 => (x"c1",x"9c",x"ff",x"ff"),
   298 => (x"c1",x"34",x"ca",x"84"),
   299 => (x"dc",x"c2",x"87",x"e7"),
   300 => (x"49",x"bf",x"97",x"e9"),
   301 => (x"99",x"c6",x"31",x"c1"),
   302 => (x"97",x"ea",x"dc",x"c2"),
   303 => (x"b7",x"c7",x"4a",x"bf"),
   304 => (x"c2",x"b1",x"72",x"2a"),
   305 => (x"bf",x"97",x"e5",x"dc"),
   306 => (x"9d",x"cf",x"4d",x"4a"),
   307 => (x"97",x"e6",x"dc",x"c2"),
   308 => (x"9a",x"c3",x"4a",x"bf"),
   309 => (x"dc",x"c2",x"32",x"ca"),
   310 => (x"4b",x"bf",x"97",x"e7"),
   311 => (x"b2",x"73",x"33",x"c2"),
   312 => (x"97",x"e8",x"dc",x"c2"),
   313 => (x"c0",x"c3",x"4b",x"bf"),
   314 => (x"2b",x"b7",x"c6",x"9b"),
   315 => (x"81",x"c2",x"b2",x"73"),
   316 => (x"30",x"71",x"48",x"c1"),
   317 => (x"48",x"c1",x"49",x"70"),
   318 => (x"4d",x"70",x"30",x"75"),
   319 => (x"84",x"c1",x"4c",x"72"),
   320 => (x"c0",x"c8",x"94",x"71"),
   321 => (x"cc",x"06",x"ad",x"b7"),
   322 => (x"b7",x"34",x"c1",x"87"),
   323 => (x"b7",x"c0",x"c8",x"2d"),
   324 => (x"f4",x"ff",x"01",x"ad"),
   325 => (x"f0",x"48",x"74",x"87"),
   326 => (x"5e",x"0e",x"87",x"d7"),
   327 => (x"0e",x"5d",x"5c",x"5b"),
   328 => (x"e5",x"c2",x"86",x"f8"),
   329 => (x"78",x"c0",x"48",x"c6"),
   330 => (x"1e",x"fe",x"dc",x"c2"),
   331 => (x"de",x"fb",x"49",x"c0"),
   332 => (x"70",x"86",x"c4",x"87"),
   333 => (x"87",x"c5",x"05",x"98"),
   334 => (x"c0",x"c9",x"48",x"c0"),
   335 => (x"c1",x"4d",x"c0",x"87"),
   336 => (x"dd",x"f2",x"c0",x"7e"),
   337 => (x"dd",x"c2",x"49",x"bf"),
   338 => (x"c8",x"71",x"4a",x"f4"),
   339 => (x"87",x"d9",x"ec",x"4b"),
   340 => (x"c2",x"05",x"98",x"70"),
   341 => (x"c0",x"7e",x"c0",x"87"),
   342 => (x"49",x"bf",x"d9",x"f2"),
   343 => (x"4a",x"d0",x"de",x"c2"),
   344 => (x"ec",x"4b",x"c8",x"71"),
   345 => (x"98",x"70",x"87",x"c3"),
   346 => (x"c0",x"87",x"c2",x"05"),
   347 => (x"c0",x"02",x"6e",x"7e"),
   348 => (x"e4",x"c2",x"87",x"fd"),
   349 => (x"c2",x"4d",x"bf",x"c4"),
   350 => (x"bf",x"9f",x"fc",x"e4"),
   351 => (x"d6",x"c5",x"48",x"7e"),
   352 => (x"c7",x"05",x"a8",x"ea"),
   353 => (x"c4",x"e4",x"c2",x"87"),
   354 => (x"87",x"ce",x"4d",x"bf"),
   355 => (x"e9",x"ca",x"48",x"6e"),
   356 => (x"c5",x"02",x"a8",x"d5"),
   357 => (x"c7",x"48",x"c0",x"87"),
   358 => (x"dc",x"c2",x"87",x"e3"),
   359 => (x"49",x"75",x"1e",x"fe"),
   360 => (x"c4",x"87",x"ec",x"f9"),
   361 => (x"05",x"98",x"70",x"86"),
   362 => (x"48",x"c0",x"87",x"c5"),
   363 => (x"c0",x"87",x"ce",x"c7"),
   364 => (x"49",x"bf",x"d9",x"f2"),
   365 => (x"4a",x"d0",x"de",x"c2"),
   366 => (x"ea",x"4b",x"c8",x"71"),
   367 => (x"98",x"70",x"87",x"eb"),
   368 => (x"c2",x"87",x"c8",x"05"),
   369 => (x"c1",x"48",x"c6",x"e5"),
   370 => (x"c0",x"87",x"da",x"78"),
   371 => (x"49",x"bf",x"dd",x"f2"),
   372 => (x"4a",x"f4",x"dd",x"c2"),
   373 => (x"ea",x"4b",x"c8",x"71"),
   374 => (x"98",x"70",x"87",x"cf"),
   375 => (x"87",x"c5",x"c0",x"02"),
   376 => (x"d8",x"c6",x"48",x"c0"),
   377 => (x"fc",x"e4",x"c2",x"87"),
   378 => (x"c1",x"49",x"bf",x"97"),
   379 => (x"c0",x"05",x"a9",x"d5"),
   380 => (x"e4",x"c2",x"87",x"cd"),
   381 => (x"49",x"bf",x"97",x"fd"),
   382 => (x"02",x"a9",x"ea",x"c2"),
   383 => (x"c0",x"87",x"c5",x"c0"),
   384 => (x"87",x"f9",x"c5",x"48"),
   385 => (x"97",x"fe",x"dc",x"c2"),
   386 => (x"c3",x"48",x"7e",x"bf"),
   387 => (x"c0",x"02",x"a8",x"e9"),
   388 => (x"48",x"6e",x"87",x"ce"),
   389 => (x"02",x"a8",x"eb",x"c3"),
   390 => (x"c0",x"87",x"c5",x"c0"),
   391 => (x"87",x"dd",x"c5",x"48"),
   392 => (x"97",x"c9",x"dd",x"c2"),
   393 => (x"05",x"99",x"49",x"bf"),
   394 => (x"c2",x"87",x"cc",x"c0"),
   395 => (x"bf",x"97",x"ca",x"dd"),
   396 => (x"02",x"a9",x"c2",x"49"),
   397 => (x"c0",x"87",x"c5",x"c0"),
   398 => (x"87",x"c1",x"c5",x"48"),
   399 => (x"97",x"cb",x"dd",x"c2"),
   400 => (x"e5",x"c2",x"48",x"bf"),
   401 => (x"4c",x"70",x"58",x"c2"),
   402 => (x"c2",x"88",x"c1",x"48"),
   403 => (x"c2",x"58",x"c6",x"e5"),
   404 => (x"bf",x"97",x"cc",x"dd"),
   405 => (x"c2",x"81",x"75",x"49"),
   406 => (x"bf",x"97",x"cd",x"dd"),
   407 => (x"72",x"32",x"c8",x"4a"),
   408 => (x"e9",x"c2",x"7e",x"a1"),
   409 => (x"78",x"6e",x"48",x"d3"),
   410 => (x"97",x"ce",x"dd",x"c2"),
   411 => (x"a6",x"c8",x"48",x"bf"),
   412 => (x"c6",x"e5",x"c2",x"58"),
   413 => (x"cf",x"c2",x"02",x"bf"),
   414 => (x"d9",x"f2",x"c0",x"87"),
   415 => (x"de",x"c2",x"49",x"bf"),
   416 => (x"c8",x"71",x"4a",x"d0"),
   417 => (x"87",x"e1",x"e7",x"4b"),
   418 => (x"c0",x"02",x"98",x"70"),
   419 => (x"48",x"c0",x"87",x"c5"),
   420 => (x"c2",x"87",x"ea",x"c3"),
   421 => (x"4c",x"bf",x"fe",x"e4"),
   422 => (x"5c",x"e7",x"e9",x"c2"),
   423 => (x"97",x"e3",x"dd",x"c2"),
   424 => (x"31",x"c8",x"49",x"bf"),
   425 => (x"97",x"e2",x"dd",x"c2"),
   426 => (x"49",x"a1",x"4a",x"bf"),
   427 => (x"97",x"e4",x"dd",x"c2"),
   428 => (x"32",x"d0",x"4a",x"bf"),
   429 => (x"c2",x"49",x"a1",x"72"),
   430 => (x"bf",x"97",x"e5",x"dd"),
   431 => (x"72",x"32",x"d8",x"4a"),
   432 => (x"66",x"c4",x"49",x"a1"),
   433 => (x"d3",x"e9",x"c2",x"91"),
   434 => (x"e9",x"c2",x"81",x"bf"),
   435 => (x"dd",x"c2",x"59",x"db"),
   436 => (x"4a",x"bf",x"97",x"eb"),
   437 => (x"dd",x"c2",x"32",x"c8"),
   438 => (x"4b",x"bf",x"97",x"ea"),
   439 => (x"dd",x"c2",x"4a",x"a2"),
   440 => (x"4b",x"bf",x"97",x"ec"),
   441 => (x"a2",x"73",x"33",x"d0"),
   442 => (x"ed",x"dd",x"c2",x"4a"),
   443 => (x"cf",x"4b",x"bf",x"97"),
   444 => (x"73",x"33",x"d8",x"9b"),
   445 => (x"e9",x"c2",x"4a",x"a2"),
   446 => (x"8a",x"c2",x"5a",x"df"),
   447 => (x"e9",x"c2",x"92",x"74"),
   448 => (x"a1",x"72",x"48",x"df"),
   449 => (x"87",x"c1",x"c1",x"78"),
   450 => (x"97",x"d0",x"dd",x"c2"),
   451 => (x"31",x"c8",x"49",x"bf"),
   452 => (x"97",x"cf",x"dd",x"c2"),
   453 => (x"49",x"a1",x"4a",x"bf"),
   454 => (x"ff",x"c7",x"31",x"c5"),
   455 => (x"c2",x"29",x"c9",x"81"),
   456 => (x"c2",x"59",x"e7",x"e9"),
   457 => (x"bf",x"97",x"d5",x"dd"),
   458 => (x"c2",x"32",x"c8",x"4a"),
   459 => (x"bf",x"97",x"d4",x"dd"),
   460 => (x"c4",x"4a",x"a2",x"4b"),
   461 => (x"82",x"6e",x"92",x"66"),
   462 => (x"5a",x"e3",x"e9",x"c2"),
   463 => (x"48",x"db",x"e9",x"c2"),
   464 => (x"e9",x"c2",x"78",x"c0"),
   465 => (x"a1",x"72",x"48",x"d7"),
   466 => (x"e7",x"e9",x"c2",x"78"),
   467 => (x"db",x"e9",x"c2",x"48"),
   468 => (x"e9",x"c2",x"78",x"bf"),
   469 => (x"e9",x"c2",x"48",x"eb"),
   470 => (x"c2",x"78",x"bf",x"df"),
   471 => (x"02",x"bf",x"c6",x"e5"),
   472 => (x"74",x"87",x"c9",x"c0"),
   473 => (x"70",x"30",x"c4",x"48"),
   474 => (x"87",x"c9",x"c0",x"7e"),
   475 => (x"bf",x"e3",x"e9",x"c2"),
   476 => (x"70",x"30",x"c4",x"48"),
   477 => (x"ca",x"e5",x"c2",x"7e"),
   478 => (x"c1",x"78",x"6e",x"48"),
   479 => (x"26",x"8e",x"f8",x"48"),
   480 => (x"26",x"4c",x"26",x"4d"),
   481 => (x"0e",x"4f",x"26",x"4b"),
   482 => (x"5d",x"5c",x"5b",x"5e"),
   483 => (x"c2",x"4a",x"71",x"0e"),
   484 => (x"02",x"bf",x"c6",x"e5"),
   485 => (x"4b",x"72",x"87",x"cb"),
   486 => (x"4d",x"72",x"2b",x"c7"),
   487 => (x"c9",x"9d",x"ff",x"c1"),
   488 => (x"c8",x"4b",x"72",x"87"),
   489 => (x"c3",x"4d",x"72",x"2b"),
   490 => (x"e9",x"c2",x"9d",x"ff"),
   491 => (x"c0",x"83",x"bf",x"d3"),
   492 => (x"ab",x"bf",x"d5",x"f2"),
   493 => (x"c0",x"87",x"d9",x"02"),
   494 => (x"c2",x"5b",x"d9",x"f2"),
   495 => (x"73",x"1e",x"fe",x"dc"),
   496 => (x"87",x"cb",x"f1",x"49"),
   497 => (x"98",x"70",x"86",x"c4"),
   498 => (x"c0",x"87",x"c5",x"05"),
   499 => (x"87",x"e6",x"c0",x"48"),
   500 => (x"bf",x"c6",x"e5",x"c2"),
   501 => (x"75",x"87",x"d2",x"02"),
   502 => (x"c2",x"91",x"c4",x"49"),
   503 => (x"69",x"81",x"fe",x"dc"),
   504 => (x"ff",x"ff",x"cf",x"4c"),
   505 => (x"cb",x"9c",x"ff",x"ff"),
   506 => (x"c2",x"49",x"75",x"87"),
   507 => (x"fe",x"dc",x"c2",x"91"),
   508 => (x"4c",x"69",x"9f",x"81"),
   509 => (x"c6",x"fe",x"48",x"74"),
   510 => (x"5b",x"5e",x"0e",x"87"),
   511 => (x"f8",x"0e",x"5d",x"5c"),
   512 => (x"9c",x"4c",x"71",x"86"),
   513 => (x"c0",x"87",x"c5",x"05"),
   514 => (x"87",x"c0",x"c3",x"48"),
   515 => (x"48",x"7e",x"a4",x"c8"),
   516 => (x"66",x"d8",x"78",x"c0"),
   517 => (x"d8",x"87",x"c7",x"02"),
   518 => (x"05",x"bf",x"97",x"66"),
   519 => (x"48",x"c0",x"87",x"c5"),
   520 => (x"c0",x"87",x"e9",x"c2"),
   521 => (x"49",x"49",x"c1",x"1e"),
   522 => (x"c4",x"87",x"d3",x"ca"),
   523 => (x"9d",x"4d",x"70",x"86"),
   524 => (x"87",x"c2",x"c1",x"02"),
   525 => (x"4a",x"ce",x"e5",x"c2"),
   526 => (x"e0",x"49",x"66",x"d8"),
   527 => (x"98",x"70",x"87",x"d0"),
   528 => (x"87",x"f2",x"c0",x"02"),
   529 => (x"66",x"d8",x"4a",x"75"),
   530 => (x"e0",x"4b",x"cb",x"49"),
   531 => (x"98",x"70",x"87",x"f5"),
   532 => (x"87",x"e2",x"c0",x"02"),
   533 => (x"9d",x"75",x"1e",x"c0"),
   534 => (x"c8",x"87",x"c7",x"02"),
   535 => (x"78",x"c0",x"48",x"a6"),
   536 => (x"a6",x"c8",x"87",x"c5"),
   537 => (x"c8",x"78",x"c1",x"48"),
   538 => (x"d1",x"c9",x"49",x"66"),
   539 => (x"70",x"86",x"c4",x"87"),
   540 => (x"fe",x"05",x"9d",x"4d"),
   541 => (x"9d",x"75",x"87",x"fe"),
   542 => (x"87",x"ce",x"c1",x"02"),
   543 => (x"6e",x"49",x"a5",x"dc"),
   544 => (x"da",x"78",x"69",x"48"),
   545 => (x"a6",x"c4",x"49",x"a5"),
   546 => (x"78",x"a4",x"c4",x"48"),
   547 => (x"c4",x"48",x"69",x"9f"),
   548 => (x"c2",x"78",x"08",x"66"),
   549 => (x"02",x"bf",x"c6",x"e5"),
   550 => (x"a5",x"d4",x"87",x"d2"),
   551 => (x"49",x"69",x"9f",x"49"),
   552 => (x"99",x"ff",x"ff",x"c0"),
   553 => (x"30",x"d0",x"48",x"71"),
   554 => (x"87",x"c2",x"7e",x"70"),
   555 => (x"48",x"6e",x"7e",x"c0"),
   556 => (x"80",x"bf",x"66",x"c4"),
   557 => (x"78",x"08",x"66",x"c4"),
   558 => (x"a4",x"cc",x"7c",x"c0"),
   559 => (x"bf",x"66",x"c4",x"49"),
   560 => (x"49",x"a4",x"d0",x"79"),
   561 => (x"48",x"c1",x"79",x"c0"),
   562 => (x"48",x"c0",x"87",x"c2"),
   563 => (x"ee",x"fa",x"8e",x"f8"),
   564 => (x"5b",x"5e",x"0e",x"87"),
   565 => (x"4c",x"71",x"0e",x"5c"),
   566 => (x"cb",x"c1",x"02",x"9c"),
   567 => (x"49",x"a4",x"c8",x"87"),
   568 => (x"c3",x"c1",x"02",x"69"),
   569 => (x"cc",x"49",x"6c",x"87"),
   570 => (x"80",x"71",x"48",x"66"),
   571 => (x"70",x"58",x"a6",x"d0"),
   572 => (x"c2",x"e5",x"c2",x"b9"),
   573 => (x"ba",x"ff",x"4a",x"bf"),
   574 => (x"99",x"71",x"99",x"72"),
   575 => (x"87",x"e5",x"c0",x"02"),
   576 => (x"6b",x"4b",x"a4",x"c4"),
   577 => (x"87",x"ff",x"f9",x"49"),
   578 => (x"e4",x"c2",x"7b",x"70"),
   579 => (x"6c",x"49",x"bf",x"fe"),
   580 => (x"cc",x"7c",x"71",x"81"),
   581 => (x"e5",x"c2",x"b9",x"66"),
   582 => (x"ff",x"4a",x"bf",x"c2"),
   583 => (x"71",x"99",x"72",x"ba"),
   584 => (x"db",x"ff",x"05",x"99"),
   585 => (x"7c",x"66",x"cc",x"87"),
   586 => (x"1e",x"87",x"d6",x"f9"),
   587 => (x"4b",x"71",x"1e",x"73"),
   588 => (x"87",x"c7",x"02",x"9b"),
   589 => (x"69",x"49",x"a3",x"c8"),
   590 => (x"c0",x"87",x"c5",x"05"),
   591 => (x"87",x"f6",x"c0",x"48"),
   592 => (x"bf",x"d7",x"e9",x"c2"),
   593 => (x"4a",x"a3",x"c4",x"49"),
   594 => (x"8a",x"c2",x"4a",x"6a"),
   595 => (x"bf",x"fe",x"e4",x"c2"),
   596 => (x"49",x"a1",x"72",x"92"),
   597 => (x"bf",x"c2",x"e5",x"c2"),
   598 => (x"72",x"9a",x"6b",x"4a"),
   599 => (x"f2",x"c0",x"49",x"a1"),
   600 => (x"66",x"c8",x"59",x"d9"),
   601 => (x"e6",x"ea",x"71",x"1e"),
   602 => (x"70",x"86",x"c4",x"87"),
   603 => (x"87",x"c4",x"05",x"98"),
   604 => (x"87",x"c2",x"48",x"c0"),
   605 => (x"ca",x"f8",x"48",x"c1"),
   606 => (x"1e",x"73",x"1e",x"87"),
   607 => (x"02",x"9b",x"4b",x"71"),
   608 => (x"a3",x"c8",x"87",x"c7"),
   609 => (x"c5",x"05",x"69",x"49"),
   610 => (x"c0",x"48",x"c0",x"87"),
   611 => (x"e9",x"c2",x"87",x"f6"),
   612 => (x"c4",x"49",x"bf",x"d7"),
   613 => (x"4a",x"6a",x"4a",x"a3"),
   614 => (x"e4",x"c2",x"8a",x"c2"),
   615 => (x"72",x"92",x"bf",x"fe"),
   616 => (x"e5",x"c2",x"49",x"a1"),
   617 => (x"6b",x"4a",x"bf",x"c2"),
   618 => (x"49",x"a1",x"72",x"9a"),
   619 => (x"59",x"d9",x"f2",x"c0"),
   620 => (x"71",x"1e",x"66",x"c8"),
   621 => (x"c4",x"87",x"d1",x"e6"),
   622 => (x"05",x"98",x"70",x"86"),
   623 => (x"48",x"c0",x"87",x"c4"),
   624 => (x"48",x"c1",x"87",x"c2"),
   625 => (x"0e",x"87",x"fc",x"f6"),
   626 => (x"5d",x"5c",x"5b",x"5e"),
   627 => (x"4b",x"71",x"1e",x"0e"),
   628 => (x"73",x"4d",x"66",x"d4"),
   629 => (x"cc",x"c1",x"02",x"9b"),
   630 => (x"49",x"a3",x"c8",x"87"),
   631 => (x"c4",x"c1",x"02",x"69"),
   632 => (x"4c",x"a3",x"d0",x"87"),
   633 => (x"bf",x"c2",x"e5",x"c2"),
   634 => (x"6c",x"b9",x"ff",x"49"),
   635 => (x"d4",x"7e",x"99",x"4a"),
   636 => (x"cd",x"06",x"a9",x"66"),
   637 => (x"7c",x"7b",x"c0",x"87"),
   638 => (x"c4",x"4a",x"a3",x"cc"),
   639 => (x"79",x"6a",x"49",x"a3"),
   640 => (x"49",x"72",x"87",x"ca"),
   641 => (x"d4",x"99",x"c0",x"f8"),
   642 => (x"8d",x"71",x"4d",x"66"),
   643 => (x"29",x"c9",x"49",x"75"),
   644 => (x"49",x"73",x"1e",x"71"),
   645 => (x"c2",x"87",x"fa",x"fa"),
   646 => (x"73",x"1e",x"fe",x"dc"),
   647 => (x"87",x"cb",x"fc",x"49"),
   648 => (x"66",x"d4",x"86",x"c8"),
   649 => (x"d6",x"f5",x"26",x"7c"),
   650 => (x"1e",x"73",x"1e",x"87"),
   651 => (x"02",x"9b",x"4b",x"71"),
   652 => (x"c2",x"87",x"e4",x"c0"),
   653 => (x"73",x"5b",x"eb",x"e9"),
   654 => (x"c2",x"8a",x"c2",x"4a"),
   655 => (x"49",x"bf",x"fe",x"e4"),
   656 => (x"d7",x"e9",x"c2",x"92"),
   657 => (x"80",x"72",x"48",x"bf"),
   658 => (x"58",x"ef",x"e9",x"c2"),
   659 => (x"30",x"c4",x"48",x"71"),
   660 => (x"58",x"ce",x"e5",x"c2"),
   661 => (x"c2",x"87",x"ed",x"c0"),
   662 => (x"c2",x"48",x"e7",x"e9"),
   663 => (x"78",x"bf",x"db",x"e9"),
   664 => (x"48",x"eb",x"e9",x"c2"),
   665 => (x"bf",x"df",x"e9",x"c2"),
   666 => (x"c6",x"e5",x"c2",x"78"),
   667 => (x"87",x"c9",x"02",x"bf"),
   668 => (x"bf",x"fe",x"e4",x"c2"),
   669 => (x"c7",x"31",x"c4",x"49"),
   670 => (x"e3",x"e9",x"c2",x"87"),
   671 => (x"31",x"c4",x"49",x"bf"),
   672 => (x"59",x"ce",x"e5",x"c2"),
   673 => (x"0e",x"87",x"fc",x"f3"),
   674 => (x"0e",x"5c",x"5b",x"5e"),
   675 => (x"4b",x"c0",x"4a",x"71"),
   676 => (x"c0",x"02",x"9a",x"72"),
   677 => (x"a2",x"da",x"87",x"e0"),
   678 => (x"4b",x"69",x"9f",x"49"),
   679 => (x"bf",x"c6",x"e5",x"c2"),
   680 => (x"d4",x"87",x"cf",x"02"),
   681 => (x"69",x"9f",x"49",x"a2"),
   682 => (x"ff",x"c0",x"4c",x"49"),
   683 => (x"34",x"d0",x"9c",x"ff"),
   684 => (x"4c",x"c0",x"87",x"c2"),
   685 => (x"49",x"73",x"b3",x"74"),
   686 => (x"f3",x"87",x"ee",x"fd"),
   687 => (x"5e",x"0e",x"87",x"c3"),
   688 => (x"0e",x"5d",x"5c",x"5b"),
   689 => (x"4a",x"71",x"86",x"f4"),
   690 => (x"9a",x"72",x"7e",x"c0"),
   691 => (x"c2",x"87",x"d8",x"02"),
   692 => (x"c0",x"48",x"fa",x"dc"),
   693 => (x"f2",x"dc",x"c2",x"78"),
   694 => (x"eb",x"e9",x"c2",x"48"),
   695 => (x"dc",x"c2",x"78",x"bf"),
   696 => (x"e9",x"c2",x"48",x"f6"),
   697 => (x"c2",x"78",x"bf",x"e7"),
   698 => (x"c0",x"48",x"db",x"e5"),
   699 => (x"ca",x"e5",x"c2",x"50"),
   700 => (x"dc",x"c2",x"49",x"bf"),
   701 => (x"71",x"4a",x"bf",x"fa"),
   702 => (x"c9",x"c4",x"03",x"aa"),
   703 => (x"cf",x"49",x"72",x"87"),
   704 => (x"e9",x"c0",x"05",x"99"),
   705 => (x"d5",x"f2",x"c0",x"87"),
   706 => (x"f2",x"dc",x"c2",x"48"),
   707 => (x"dc",x"c2",x"78",x"bf"),
   708 => (x"dc",x"c2",x"1e",x"fe"),
   709 => (x"c2",x"49",x"bf",x"f2"),
   710 => (x"c1",x"48",x"f2",x"dc"),
   711 => (x"e3",x"71",x"78",x"a1"),
   712 => (x"86",x"c4",x"87",x"ed"),
   713 => (x"48",x"d1",x"f2",x"c0"),
   714 => (x"78",x"fe",x"dc",x"c2"),
   715 => (x"f2",x"c0",x"87",x"cc"),
   716 => (x"c0",x"48",x"bf",x"d1"),
   717 => (x"f2",x"c0",x"80",x"e0"),
   718 => (x"dc",x"c2",x"58",x"d5"),
   719 => (x"c1",x"48",x"bf",x"fa"),
   720 => (x"fe",x"dc",x"c2",x"80"),
   721 => (x"0c",x"91",x"27",x"58"),
   722 => (x"97",x"bf",x"00",x"00"),
   723 => (x"02",x"9d",x"4d",x"bf"),
   724 => (x"c3",x"87",x"e3",x"c2"),
   725 => (x"c2",x"02",x"ad",x"e5"),
   726 => (x"f2",x"c0",x"87",x"dc"),
   727 => (x"cb",x"4b",x"bf",x"d1"),
   728 => (x"4c",x"11",x"49",x"a3"),
   729 => (x"c1",x"05",x"ac",x"cf"),
   730 => (x"49",x"75",x"87",x"d2"),
   731 => (x"89",x"c1",x"99",x"df"),
   732 => (x"e5",x"c2",x"91",x"cd"),
   733 => (x"a3",x"c1",x"81",x"ce"),
   734 => (x"c3",x"51",x"12",x"4a"),
   735 => (x"51",x"12",x"4a",x"a3"),
   736 => (x"12",x"4a",x"a3",x"c5"),
   737 => (x"4a",x"a3",x"c7",x"51"),
   738 => (x"a3",x"c9",x"51",x"12"),
   739 => (x"ce",x"51",x"12",x"4a"),
   740 => (x"51",x"12",x"4a",x"a3"),
   741 => (x"12",x"4a",x"a3",x"d0"),
   742 => (x"4a",x"a3",x"d2",x"51"),
   743 => (x"a3",x"d4",x"51",x"12"),
   744 => (x"d6",x"51",x"12",x"4a"),
   745 => (x"51",x"12",x"4a",x"a3"),
   746 => (x"12",x"4a",x"a3",x"d8"),
   747 => (x"4a",x"a3",x"dc",x"51"),
   748 => (x"a3",x"de",x"51",x"12"),
   749 => (x"c1",x"51",x"12",x"4a"),
   750 => (x"87",x"fa",x"c0",x"7e"),
   751 => (x"99",x"c8",x"49",x"74"),
   752 => (x"87",x"eb",x"c0",x"05"),
   753 => (x"99",x"d0",x"49",x"74"),
   754 => (x"dc",x"87",x"d1",x"05"),
   755 => (x"cb",x"c0",x"02",x"66"),
   756 => (x"dc",x"49",x"73",x"87"),
   757 => (x"98",x"70",x"0f",x"66"),
   758 => (x"87",x"d3",x"c0",x"02"),
   759 => (x"c6",x"c0",x"05",x"6e"),
   760 => (x"ce",x"e5",x"c2",x"87"),
   761 => (x"c0",x"50",x"c0",x"48"),
   762 => (x"48",x"bf",x"d1",x"f2"),
   763 => (x"c2",x"87",x"dd",x"c2"),
   764 => (x"c0",x"48",x"db",x"e5"),
   765 => (x"e5",x"c2",x"7e",x"50"),
   766 => (x"c2",x"49",x"bf",x"ca"),
   767 => (x"4a",x"bf",x"fa",x"dc"),
   768 => (x"fb",x"04",x"aa",x"71"),
   769 => (x"e9",x"c2",x"87",x"f7"),
   770 => (x"c0",x"05",x"bf",x"eb"),
   771 => (x"e5",x"c2",x"87",x"c8"),
   772 => (x"c1",x"02",x"bf",x"c6"),
   773 => (x"dc",x"c2",x"87",x"f4"),
   774 => (x"ed",x"49",x"bf",x"f6"),
   775 => (x"dc",x"c2",x"87",x"e9"),
   776 => (x"a6",x"c4",x"58",x"fa"),
   777 => (x"f6",x"dc",x"c2",x"48"),
   778 => (x"e5",x"c2",x"78",x"bf"),
   779 => (x"c0",x"02",x"bf",x"c6"),
   780 => (x"66",x"c4",x"87",x"d8"),
   781 => (x"ff",x"ff",x"cf",x"49"),
   782 => (x"a9",x"99",x"f8",x"ff"),
   783 => (x"87",x"c5",x"c0",x"02"),
   784 => (x"e1",x"c0",x"4c",x"c0"),
   785 => (x"c0",x"4c",x"c1",x"87"),
   786 => (x"66",x"c4",x"87",x"dc"),
   787 => (x"f8",x"ff",x"cf",x"49"),
   788 => (x"c0",x"02",x"a9",x"99"),
   789 => (x"a6",x"c8",x"87",x"c8"),
   790 => (x"c0",x"78",x"c0",x"48"),
   791 => (x"a6",x"c8",x"87",x"c5"),
   792 => (x"c8",x"78",x"c1",x"48"),
   793 => (x"9c",x"74",x"4c",x"66"),
   794 => (x"87",x"de",x"c0",x"05"),
   795 => (x"c2",x"49",x"66",x"c4"),
   796 => (x"fe",x"e4",x"c2",x"89"),
   797 => (x"e9",x"c2",x"91",x"bf"),
   798 => (x"71",x"48",x"bf",x"d7"),
   799 => (x"f6",x"dc",x"c2",x"80"),
   800 => (x"fa",x"dc",x"c2",x"58"),
   801 => (x"f9",x"78",x"c0",x"48"),
   802 => (x"48",x"c0",x"87",x"e3"),
   803 => (x"ee",x"eb",x"8e",x"f4"),
   804 => (x"00",x"00",x"00",x"87"),
   805 => (x"ff",x"ff",x"ff",x"00"),
   806 => (x"00",x"0c",x"a1",x"ff"),
   807 => (x"00",x"0c",x"aa",x"00"),
   808 => (x"54",x"41",x"46",x"00"),
   809 => (x"20",x"20",x"32",x"33"),
   810 => (x"41",x"46",x"00",x"20"),
   811 => (x"20",x"36",x"31",x"54"),
   812 => (x"1e",x"00",x"20",x"20"),
   813 => (x"c3",x"48",x"d4",x"ff"),
   814 => (x"48",x"68",x"78",x"ff"),
   815 => (x"ff",x"1e",x"4f",x"26"),
   816 => (x"ff",x"c3",x"48",x"d4"),
   817 => (x"48",x"d0",x"ff",x"78"),
   818 => (x"ff",x"78",x"e1",x"c0"),
   819 => (x"78",x"d4",x"48",x"d4"),
   820 => (x"48",x"ef",x"e9",x"c2"),
   821 => (x"50",x"bf",x"d4",x"ff"),
   822 => (x"ff",x"1e",x"4f",x"26"),
   823 => (x"e0",x"c0",x"48",x"d0"),
   824 => (x"1e",x"4f",x"26",x"78"),
   825 => (x"70",x"87",x"cc",x"ff"),
   826 => (x"c6",x"02",x"99",x"49"),
   827 => (x"a9",x"fb",x"c0",x"87"),
   828 => (x"71",x"87",x"f1",x"05"),
   829 => (x"0e",x"4f",x"26",x"48"),
   830 => (x"0e",x"5c",x"5b",x"5e"),
   831 => (x"4c",x"c0",x"4b",x"71"),
   832 => (x"70",x"87",x"f0",x"fe"),
   833 => (x"c0",x"02",x"99",x"49"),
   834 => (x"ec",x"c0",x"87",x"f9"),
   835 => (x"f2",x"c0",x"02",x"a9"),
   836 => (x"a9",x"fb",x"c0",x"87"),
   837 => (x"87",x"eb",x"c0",x"02"),
   838 => (x"ac",x"b7",x"66",x"cc"),
   839 => (x"d0",x"87",x"c7",x"03"),
   840 => (x"87",x"c2",x"02",x"66"),
   841 => (x"99",x"71",x"53",x"71"),
   842 => (x"c1",x"87",x"c2",x"02"),
   843 => (x"87",x"c3",x"fe",x"84"),
   844 => (x"02",x"99",x"49",x"70"),
   845 => (x"ec",x"c0",x"87",x"cd"),
   846 => (x"87",x"c7",x"02",x"a9"),
   847 => (x"05",x"a9",x"fb",x"c0"),
   848 => (x"d0",x"87",x"d5",x"ff"),
   849 => (x"87",x"c3",x"02",x"66"),
   850 => (x"c0",x"7b",x"97",x"c0"),
   851 => (x"c4",x"05",x"a9",x"ec"),
   852 => (x"c5",x"4a",x"74",x"87"),
   853 => (x"c0",x"4a",x"74",x"87"),
   854 => (x"48",x"72",x"8a",x"0a"),
   855 => (x"4d",x"26",x"87",x"c2"),
   856 => (x"4b",x"26",x"4c",x"26"),
   857 => (x"fd",x"1e",x"4f",x"26"),
   858 => (x"49",x"70",x"87",x"c9"),
   859 => (x"aa",x"f0",x"c0",x"4a"),
   860 => (x"c0",x"87",x"c9",x"04"),
   861 => (x"c3",x"01",x"aa",x"f9"),
   862 => (x"8a",x"f0",x"c0",x"87"),
   863 => (x"04",x"aa",x"c1",x"c1"),
   864 => (x"da",x"c1",x"87",x"c9"),
   865 => (x"87",x"c3",x"01",x"aa"),
   866 => (x"72",x"8a",x"f7",x"c0"),
   867 => (x"0e",x"4f",x"26",x"48"),
   868 => (x"0e",x"5c",x"5b",x"5e"),
   869 => (x"d4",x"ff",x"4a",x"71"),
   870 => (x"c0",x"49",x"72",x"4b"),
   871 => (x"4c",x"70",x"87",x"e7"),
   872 => (x"87",x"c2",x"02",x"9c"),
   873 => (x"d0",x"ff",x"8c",x"c1"),
   874 => (x"c1",x"78",x"c5",x"48"),
   875 => (x"49",x"74",x"7b",x"d5"),
   876 => (x"e3",x"c1",x"31",x"c6"),
   877 => (x"4a",x"bf",x"97",x"dc"),
   878 => (x"70",x"b0",x"71",x"48"),
   879 => (x"48",x"d0",x"ff",x"7b"),
   880 => (x"db",x"fe",x"78",x"c4"),
   881 => (x"5b",x"5e",x"0e",x"87"),
   882 => (x"f8",x"0e",x"5d",x"5c"),
   883 => (x"c0",x"4c",x"71",x"86"),
   884 => (x"87",x"ea",x"fb",x"7e"),
   885 => (x"f9",x"c0",x"4b",x"c0"),
   886 => (x"49",x"bf",x"97",x"f2"),
   887 => (x"cf",x"04",x"a9",x"c0"),
   888 => (x"87",x"ff",x"fb",x"87"),
   889 => (x"f9",x"c0",x"83",x"c1"),
   890 => (x"49",x"bf",x"97",x"f2"),
   891 => (x"87",x"f1",x"06",x"ab"),
   892 => (x"97",x"f2",x"f9",x"c0"),
   893 => (x"87",x"cf",x"02",x"bf"),
   894 => (x"70",x"87",x"f8",x"fa"),
   895 => (x"c6",x"02",x"99",x"49"),
   896 => (x"a9",x"ec",x"c0",x"87"),
   897 => (x"c0",x"87",x"f1",x"05"),
   898 => (x"87",x"e7",x"fa",x"4b"),
   899 => (x"e2",x"fa",x"4d",x"70"),
   900 => (x"58",x"a6",x"c8",x"87"),
   901 => (x"70",x"87",x"dc",x"fa"),
   902 => (x"c8",x"83",x"c1",x"4a"),
   903 => (x"69",x"97",x"49",x"a4"),
   904 => (x"c7",x"02",x"ad",x"49"),
   905 => (x"ad",x"ff",x"c0",x"87"),
   906 => (x"87",x"e7",x"c0",x"05"),
   907 => (x"97",x"49",x"a4",x"c9"),
   908 => (x"66",x"c4",x"49",x"69"),
   909 => (x"87",x"c7",x"02",x"a9"),
   910 => (x"a8",x"ff",x"c0",x"48"),
   911 => (x"ca",x"87",x"d4",x"05"),
   912 => (x"69",x"97",x"49",x"a4"),
   913 => (x"c6",x"02",x"aa",x"49"),
   914 => (x"aa",x"ff",x"c0",x"87"),
   915 => (x"c1",x"87",x"c4",x"05"),
   916 => (x"c0",x"87",x"d0",x"7e"),
   917 => (x"c6",x"02",x"ad",x"ec"),
   918 => (x"ad",x"fb",x"c0",x"87"),
   919 => (x"c0",x"87",x"c4",x"05"),
   920 => (x"6e",x"7e",x"c1",x"4b"),
   921 => (x"87",x"e1",x"fe",x"02"),
   922 => (x"73",x"87",x"ef",x"f9"),
   923 => (x"fb",x"8e",x"f8",x"48"),
   924 => (x"0e",x"00",x"87",x"ec"),
   925 => (x"5d",x"5c",x"5b",x"5e"),
   926 => (x"71",x"86",x"f8",x"0e"),
   927 => (x"4b",x"d4",x"ff",x"4d"),
   928 => (x"e9",x"c2",x"1e",x"75"),
   929 => (x"f0",x"e5",x"49",x"f4"),
   930 => (x"70",x"86",x"c4",x"87"),
   931 => (x"ca",x"c4",x"02",x"98"),
   932 => (x"48",x"a6",x"c4",x"87"),
   933 => (x"bf",x"de",x"e3",x"c1"),
   934 => (x"fb",x"49",x"75",x"78"),
   935 => (x"d0",x"ff",x"87",x"f1"),
   936 => (x"c1",x"78",x"c5",x"48"),
   937 => (x"4a",x"c0",x"7b",x"d6"),
   938 => (x"11",x"49",x"a2",x"75"),
   939 => (x"cb",x"82",x"c1",x"7b"),
   940 => (x"f3",x"04",x"aa",x"b7"),
   941 => (x"c3",x"4a",x"cc",x"87"),
   942 => (x"82",x"c1",x"7b",x"ff"),
   943 => (x"aa",x"b7",x"e0",x"c0"),
   944 => (x"ff",x"87",x"f4",x"04"),
   945 => (x"78",x"c4",x"48",x"d0"),
   946 => (x"c5",x"7b",x"ff",x"c3"),
   947 => (x"7b",x"d3",x"c1",x"78"),
   948 => (x"78",x"c4",x"7b",x"c1"),
   949 => (x"b7",x"c0",x"48",x"66"),
   950 => (x"ee",x"c2",x"06",x"a8"),
   951 => (x"fc",x"e9",x"c2",x"87"),
   952 => (x"66",x"c4",x"4c",x"bf"),
   953 => (x"c8",x"88",x"74",x"48"),
   954 => (x"9c",x"74",x"58",x"a6"),
   955 => (x"87",x"f7",x"c1",x"02"),
   956 => (x"7e",x"fe",x"dc",x"c2"),
   957 => (x"8c",x"4d",x"c0",x"c8"),
   958 => (x"03",x"ac",x"b7",x"c0"),
   959 => (x"c0",x"c8",x"87",x"c6"),
   960 => (x"4c",x"c0",x"4d",x"a4"),
   961 => (x"97",x"ef",x"e9",x"c2"),
   962 => (x"99",x"d0",x"49",x"bf"),
   963 => (x"c0",x"87",x"d0",x"02"),
   964 => (x"f4",x"e9",x"c2",x"1e"),
   965 => (x"87",x"d3",x"e8",x"49"),
   966 => (x"4a",x"70",x"86",x"c4"),
   967 => (x"c2",x"87",x"ed",x"c0"),
   968 => (x"c2",x"1e",x"fe",x"dc"),
   969 => (x"e8",x"49",x"f4",x"e9"),
   970 => (x"86",x"c4",x"87",x"c1"),
   971 => (x"d0",x"ff",x"4a",x"70"),
   972 => (x"78",x"c5",x"c8",x"48"),
   973 => (x"6e",x"7b",x"d4",x"c1"),
   974 => (x"6e",x"7b",x"bf",x"97"),
   975 => (x"70",x"80",x"c1",x"48"),
   976 => (x"05",x"8d",x"c1",x"7e"),
   977 => (x"ff",x"87",x"f0",x"ff"),
   978 => (x"78",x"c4",x"48",x"d0"),
   979 => (x"c5",x"05",x"9a",x"72"),
   980 => (x"c1",x"48",x"c0",x"87"),
   981 => (x"1e",x"c1",x"87",x"c7"),
   982 => (x"49",x"f4",x"e9",x"c2"),
   983 => (x"c4",x"87",x"f2",x"e5"),
   984 => (x"05",x"9c",x"74",x"86"),
   985 => (x"c4",x"87",x"c9",x"fe"),
   986 => (x"b7",x"c0",x"48",x"66"),
   987 => (x"87",x"d1",x"06",x"a8"),
   988 => (x"48",x"f4",x"e9",x"c2"),
   989 => (x"80",x"d0",x"78",x"c0"),
   990 => (x"80",x"f4",x"78",x"c0"),
   991 => (x"bf",x"c0",x"ea",x"c2"),
   992 => (x"48",x"66",x"c4",x"78"),
   993 => (x"01",x"a8",x"b7",x"c0"),
   994 => (x"ff",x"87",x"d2",x"fd"),
   995 => (x"78",x"c5",x"48",x"d0"),
   996 => (x"c0",x"7b",x"d3",x"c1"),
   997 => (x"c1",x"78",x"c4",x"7b"),
   998 => (x"c0",x"87",x"c2",x"48"),
   999 => (x"26",x"8e",x"f8",x"48"),
  1000 => (x"26",x"4c",x"26",x"4d"),
  1001 => (x"0e",x"4f",x"26",x"4b"),
  1002 => (x"5d",x"5c",x"5b",x"5e"),
  1003 => (x"4b",x"71",x"1e",x"0e"),
  1004 => (x"ab",x"4d",x"4c",x"c0"),
  1005 => (x"87",x"e8",x"c0",x"04"),
  1006 => (x"1e",x"c5",x"f7",x"c0"),
  1007 => (x"c4",x"02",x"9d",x"75"),
  1008 => (x"c2",x"4a",x"c0",x"87"),
  1009 => (x"72",x"4a",x"c1",x"87"),
  1010 => (x"87",x"f2",x"eb",x"49"),
  1011 => (x"7e",x"70",x"86",x"c4"),
  1012 => (x"05",x"6e",x"84",x"c1"),
  1013 => (x"4c",x"73",x"87",x"c2"),
  1014 => (x"ac",x"73",x"85",x"c1"),
  1015 => (x"87",x"d8",x"ff",x"06"),
  1016 => (x"fe",x"26",x"48",x"6e"),
  1017 => (x"5e",x"0e",x"87",x"f9"),
  1018 => (x"71",x"0e",x"5c",x"5b"),
  1019 => (x"02",x"66",x"cc",x"4b"),
  1020 => (x"c0",x"4c",x"87",x"d8"),
  1021 => (x"d8",x"02",x"8c",x"f0"),
  1022 => (x"c1",x"4a",x"74",x"87"),
  1023 => (x"87",x"d1",x"02",x"8a"),
  1024 => (x"87",x"cd",x"02",x"8a"),
  1025 => (x"87",x"c9",x"02",x"8a"),
  1026 => (x"49",x"73",x"87",x"d9"),
  1027 => (x"d2",x"87",x"e4",x"f9"),
  1028 => (x"c0",x"1e",x"74",x"87"),
  1029 => (x"d6",x"d8",x"c1",x"49"),
  1030 => (x"73",x"1e",x"74",x"87"),
  1031 => (x"ce",x"d8",x"c1",x"49"),
  1032 => (x"fd",x"86",x"c8",x"87"),
  1033 => (x"5e",x"0e",x"87",x"fb"),
  1034 => (x"0e",x"5d",x"5c",x"5b"),
  1035 => (x"49",x"4c",x"71",x"1e"),
  1036 => (x"ea",x"c2",x"91",x"de"),
  1037 => (x"85",x"71",x"4d",x"dc"),
  1038 => (x"c1",x"02",x"6d",x"97"),
  1039 => (x"ea",x"c2",x"87",x"dc"),
  1040 => (x"74",x"49",x"bf",x"c8"),
  1041 => (x"de",x"fd",x"71",x"81"),
  1042 => (x"48",x"7e",x"70",x"87"),
  1043 => (x"f2",x"c0",x"02",x"98"),
  1044 => (x"d0",x"ea",x"c2",x"87"),
  1045 => (x"cb",x"4a",x"70",x"4b"),
  1046 => (x"ca",x"c1",x"ff",x"49"),
  1047 => (x"cb",x"4b",x"74",x"87"),
  1048 => (x"f0",x"e3",x"c1",x"93"),
  1049 => (x"c1",x"83",x"c4",x"83"),
  1050 => (x"74",x"7b",x"de",x"c2"),
  1051 => (x"e5",x"c0",x"c1",x"49"),
  1052 => (x"c1",x"7b",x"75",x"87"),
  1053 => (x"bf",x"97",x"dd",x"e3"),
  1054 => (x"ea",x"c2",x"1e",x"49"),
  1055 => (x"e5",x"fd",x"49",x"d0"),
  1056 => (x"74",x"86",x"c4",x"87"),
  1057 => (x"cd",x"c0",x"c1",x"49"),
  1058 => (x"c1",x"49",x"c0",x"87"),
  1059 => (x"c2",x"87",x"ec",x"c1"),
  1060 => (x"c0",x"48",x"f0",x"e9"),
  1061 => (x"dd",x"49",x"c1",x"78"),
  1062 => (x"fc",x"26",x"87",x"fb"),
  1063 => (x"6f",x"4c",x"87",x"c1"),
  1064 => (x"6e",x"69",x"64",x"61"),
  1065 => (x"2e",x"2e",x"2e",x"67"),
  1066 => (x"1e",x"73",x"1e",x"00"),
  1067 => (x"c2",x"49",x"4a",x"71"),
  1068 => (x"81",x"bf",x"c8",x"ea"),
  1069 => (x"87",x"ef",x"fb",x"71"),
  1070 => (x"02",x"9b",x"4b",x"70"),
  1071 => (x"e7",x"49",x"87",x"c4"),
  1072 => (x"ea",x"c2",x"87",x"c5"),
  1073 => (x"78",x"c0",x"48",x"c8"),
  1074 => (x"c8",x"dd",x"49",x"c1"),
  1075 => (x"87",x"d3",x"fb",x"87"),
  1076 => (x"5c",x"5b",x"5e",x"0e"),
  1077 => (x"86",x"f4",x"0e",x"5d"),
  1078 => (x"4d",x"fe",x"dc",x"c2"),
  1079 => (x"a6",x"c4",x"4c",x"c0"),
  1080 => (x"c2",x"78",x"c0",x"48"),
  1081 => (x"48",x"bf",x"c8",x"ea"),
  1082 => (x"c1",x"06",x"a8",x"c0"),
  1083 => (x"dc",x"c2",x"87",x"c0"),
  1084 => (x"02",x"98",x"48",x"fe"),
  1085 => (x"c0",x"87",x"f7",x"c0"),
  1086 => (x"c8",x"1e",x"c5",x"f7"),
  1087 => (x"87",x"c7",x"02",x"66"),
  1088 => (x"c0",x"48",x"a6",x"c4"),
  1089 => (x"c4",x"87",x"c5",x"78"),
  1090 => (x"78",x"c1",x"48",x"a6"),
  1091 => (x"e6",x"49",x"66",x"c4"),
  1092 => (x"86",x"c4",x"87",x"ec"),
  1093 => (x"84",x"c1",x"4d",x"70"),
  1094 => (x"c1",x"48",x"66",x"c4"),
  1095 => (x"58",x"a6",x"c8",x"80"),
  1096 => (x"bf",x"c8",x"ea",x"c2"),
  1097 => (x"87",x"c6",x"03",x"ac"),
  1098 => (x"ff",x"05",x"9d",x"75"),
  1099 => (x"4c",x"c0",x"87",x"c9"),
  1100 => (x"c3",x"02",x"9d",x"75"),
  1101 => (x"f7",x"c0",x"87",x"dc"),
  1102 => (x"66",x"c8",x"1e",x"c5"),
  1103 => (x"cc",x"87",x"c7",x"02"),
  1104 => (x"78",x"c0",x"48",x"a6"),
  1105 => (x"a6",x"cc",x"87",x"c5"),
  1106 => (x"cc",x"78",x"c1",x"48"),
  1107 => (x"ed",x"e5",x"49",x"66"),
  1108 => (x"70",x"86",x"c4",x"87"),
  1109 => (x"02",x"98",x"48",x"7e"),
  1110 => (x"49",x"87",x"e4",x"c2"),
  1111 => (x"69",x"97",x"81",x"cb"),
  1112 => (x"02",x"99",x"d0",x"49"),
  1113 => (x"74",x"87",x"d4",x"c1"),
  1114 => (x"c1",x"91",x"cb",x"49"),
  1115 => (x"c1",x"81",x"f0",x"e3"),
  1116 => (x"c8",x"79",x"e9",x"c2"),
  1117 => (x"51",x"ff",x"c3",x"81"),
  1118 => (x"91",x"de",x"49",x"74"),
  1119 => (x"4d",x"dc",x"ea",x"c2"),
  1120 => (x"c1",x"c2",x"85",x"71"),
  1121 => (x"a5",x"c1",x"7d",x"97"),
  1122 => (x"51",x"e0",x"c0",x"49"),
  1123 => (x"97",x"ce",x"e5",x"c2"),
  1124 => (x"87",x"d2",x"02",x"bf"),
  1125 => (x"a5",x"c2",x"84",x"c1"),
  1126 => (x"ce",x"e5",x"c2",x"4b"),
  1127 => (x"fe",x"49",x"db",x"4a"),
  1128 => (x"c1",x"87",x"c4",x"fc"),
  1129 => (x"a5",x"cd",x"87",x"d9"),
  1130 => (x"c1",x"51",x"c0",x"49"),
  1131 => (x"4b",x"a5",x"c2",x"84"),
  1132 => (x"49",x"cb",x"4a",x"6e"),
  1133 => (x"87",x"ef",x"fb",x"fe"),
  1134 => (x"74",x"87",x"c4",x"c1"),
  1135 => (x"c1",x"91",x"cb",x"49"),
  1136 => (x"c1",x"81",x"f0",x"e3"),
  1137 => (x"c2",x"79",x"e6",x"c0"),
  1138 => (x"bf",x"97",x"ce",x"e5"),
  1139 => (x"74",x"87",x"d8",x"02"),
  1140 => (x"c1",x"91",x"de",x"49"),
  1141 => (x"dc",x"ea",x"c2",x"84"),
  1142 => (x"c2",x"83",x"71",x"4b"),
  1143 => (x"dd",x"4a",x"ce",x"e5"),
  1144 => (x"c2",x"fb",x"fe",x"49"),
  1145 => (x"74",x"87",x"d8",x"87"),
  1146 => (x"c2",x"93",x"de",x"4b"),
  1147 => (x"cb",x"83",x"dc",x"ea"),
  1148 => (x"51",x"c0",x"49",x"a3"),
  1149 => (x"6e",x"73",x"84",x"c1"),
  1150 => (x"fe",x"49",x"cb",x"4a"),
  1151 => (x"c4",x"87",x"e8",x"fa"),
  1152 => (x"80",x"c1",x"48",x"66"),
  1153 => (x"c7",x"58",x"a6",x"c8"),
  1154 => (x"c5",x"c0",x"03",x"ac"),
  1155 => (x"fc",x"05",x"6e",x"87"),
  1156 => (x"48",x"74",x"87",x"e4"),
  1157 => (x"c6",x"f6",x"8e",x"f4"),
  1158 => (x"1e",x"73",x"1e",x"87"),
  1159 => (x"cb",x"49",x"4b",x"71"),
  1160 => (x"f0",x"e3",x"c1",x"91"),
  1161 => (x"4a",x"a1",x"c8",x"81"),
  1162 => (x"48",x"dc",x"e3",x"c1"),
  1163 => (x"a1",x"c9",x"50",x"12"),
  1164 => (x"f2",x"f9",x"c0",x"4a"),
  1165 => (x"ca",x"50",x"12",x"48"),
  1166 => (x"dd",x"e3",x"c1",x"81"),
  1167 => (x"c1",x"50",x"11",x"48"),
  1168 => (x"bf",x"97",x"dd",x"e3"),
  1169 => (x"49",x"c0",x"1e",x"49"),
  1170 => (x"c2",x"87",x"db",x"f6"),
  1171 => (x"de",x"48",x"f0",x"e9"),
  1172 => (x"d6",x"49",x"c1",x"78"),
  1173 => (x"f5",x"26",x"87",x"ff"),
  1174 => (x"71",x"1e",x"87",x"c9"),
  1175 => (x"91",x"cb",x"49",x"4a"),
  1176 => (x"81",x"f0",x"e3",x"c1"),
  1177 => (x"48",x"11",x"81",x"c8"),
  1178 => (x"58",x"f4",x"e9",x"c2"),
  1179 => (x"48",x"c8",x"ea",x"c2"),
  1180 => (x"49",x"c1",x"78",x"c0"),
  1181 => (x"26",x"87",x"de",x"d6"),
  1182 => (x"49",x"c0",x"1e",x"4f"),
  1183 => (x"87",x"fb",x"f9",x"c0"),
  1184 => (x"71",x"1e",x"4f",x"26"),
  1185 => (x"87",x"d2",x"02",x"99"),
  1186 => (x"48",x"c5",x"e5",x"c1"),
  1187 => (x"80",x"f7",x"50",x"c0"),
  1188 => (x"40",x"da",x"c9",x"c1"),
  1189 => (x"78",x"e9",x"e3",x"c1"),
  1190 => (x"e5",x"c1",x"87",x"ce"),
  1191 => (x"e3",x"c1",x"48",x"c1"),
  1192 => (x"80",x"fc",x"78",x"e2"),
  1193 => (x"78",x"f9",x"c9",x"c1"),
  1194 => (x"5e",x"0e",x"4f",x"26"),
  1195 => (x"0e",x"5d",x"5c",x"5b"),
  1196 => (x"4d",x"71",x"86",x"f4"),
  1197 => (x"c1",x"91",x"cb",x"49"),
  1198 => (x"c8",x"81",x"f0",x"e3"),
  1199 => (x"a1",x"ca",x"4a",x"a1"),
  1200 => (x"48",x"a6",x"c4",x"7e"),
  1201 => (x"bf",x"f8",x"ed",x"c2"),
  1202 => (x"bf",x"97",x"6e",x"78"),
  1203 => (x"4c",x"66",x"c4",x"4b"),
  1204 => (x"48",x"12",x"2c",x"73"),
  1205 => (x"70",x"58",x"a6",x"cc"),
  1206 => (x"c9",x"84",x"c1",x"9c"),
  1207 => (x"49",x"69",x"97",x"81"),
  1208 => (x"c2",x"04",x"ac",x"b7"),
  1209 => (x"6e",x"4c",x"c0",x"87"),
  1210 => (x"c8",x"4a",x"bf",x"97"),
  1211 => (x"31",x"72",x"49",x"66"),
  1212 => (x"66",x"c4",x"b9",x"ff"),
  1213 => (x"72",x"48",x"74",x"99"),
  1214 => (x"48",x"4a",x"70",x"30"),
  1215 => (x"ed",x"c2",x"b0",x"71"),
  1216 => (x"e4",x"c0",x"58",x"fc"),
  1217 => (x"49",x"c0",x"87",x"d0"),
  1218 => (x"75",x"87",x"ca",x"d4"),
  1219 => (x"c5",x"f6",x"c0",x"49"),
  1220 => (x"f2",x"8e",x"f4",x"87"),
  1221 => (x"73",x"1e",x"87",x"c9"),
  1222 => (x"49",x"4b",x"71",x"1e"),
  1223 => (x"73",x"87",x"cb",x"fe"),
  1224 => (x"87",x"c6",x"fe",x"49"),
  1225 => (x"1e",x"87",x"fc",x"f1"),
  1226 => (x"4b",x"71",x"1e",x"73"),
  1227 => (x"02",x"4a",x"a3",x"c6"),
  1228 => (x"8a",x"c1",x"87",x"db"),
  1229 => (x"8a",x"87",x"d6",x"02"),
  1230 => (x"87",x"da",x"c1",x"02"),
  1231 => (x"fc",x"c0",x"02",x"8a"),
  1232 => (x"c0",x"02",x"8a",x"87"),
  1233 => (x"02",x"8a",x"87",x"e1"),
  1234 => (x"db",x"c1",x"87",x"cb"),
  1235 => (x"fc",x"49",x"c7",x"87"),
  1236 => (x"de",x"c1",x"87",x"c8"),
  1237 => (x"c8",x"ea",x"c2",x"87"),
  1238 => (x"cb",x"c1",x"02",x"bf"),
  1239 => (x"88",x"c1",x"48",x"87"),
  1240 => (x"58",x"cc",x"ea",x"c2"),
  1241 => (x"c2",x"87",x"c1",x"c1"),
  1242 => (x"02",x"bf",x"cc",x"ea"),
  1243 => (x"c2",x"87",x"f9",x"c0"),
  1244 => (x"48",x"bf",x"c8",x"ea"),
  1245 => (x"ea",x"c2",x"80",x"c1"),
  1246 => (x"eb",x"c0",x"58",x"cc"),
  1247 => (x"c8",x"ea",x"c2",x"87"),
  1248 => (x"89",x"c6",x"49",x"bf"),
  1249 => (x"59",x"cc",x"ea",x"c2"),
  1250 => (x"03",x"a9",x"b7",x"c0"),
  1251 => (x"ea",x"c2",x"87",x"da"),
  1252 => (x"78",x"c0",x"48",x"c8"),
  1253 => (x"ea",x"c2",x"87",x"d2"),
  1254 => (x"cb",x"02",x"bf",x"cc"),
  1255 => (x"c8",x"ea",x"c2",x"87"),
  1256 => (x"80",x"c6",x"48",x"bf"),
  1257 => (x"58",x"cc",x"ea",x"c2"),
  1258 => (x"e8",x"d1",x"49",x"c0"),
  1259 => (x"c0",x"49",x"73",x"87"),
  1260 => (x"ef",x"87",x"e3",x"f3"),
  1261 => (x"5e",x"0e",x"87",x"ed"),
  1262 => (x"0e",x"5d",x"5c",x"5b"),
  1263 => (x"dc",x"86",x"d4",x"ff"),
  1264 => (x"a6",x"c8",x"59",x"a6"),
  1265 => (x"c4",x"78",x"c0",x"48"),
  1266 => (x"66",x"c0",x"c1",x"80"),
  1267 => (x"c1",x"80",x"c4",x"78"),
  1268 => (x"c1",x"80",x"c4",x"78"),
  1269 => (x"cc",x"ea",x"c2",x"78"),
  1270 => (x"c2",x"78",x"c1",x"48"),
  1271 => (x"48",x"bf",x"f0",x"e9"),
  1272 => (x"c9",x"05",x"a8",x"de"),
  1273 => (x"87",x"e8",x"f3",x"87"),
  1274 => (x"cf",x"58",x"a6",x"cc"),
  1275 => (x"cd",x"e3",x"87",x"e6"),
  1276 => (x"87",x"ef",x"e3",x"87"),
  1277 => (x"70",x"87",x"fc",x"e2"),
  1278 => (x"ac",x"fb",x"c0",x"4c"),
  1279 => (x"87",x"fb",x"c1",x"02"),
  1280 => (x"c1",x"05",x"66",x"d8"),
  1281 => (x"fc",x"c0",x"87",x"ed"),
  1282 => (x"82",x"c4",x"4a",x"66"),
  1283 => (x"1e",x"72",x"7e",x"6a"),
  1284 => (x"48",x"c9",x"e0",x"c1"),
  1285 => (x"c8",x"49",x"66",x"c4"),
  1286 => (x"41",x"20",x"4a",x"a1"),
  1287 => (x"f9",x"05",x"aa",x"71"),
  1288 => (x"26",x"51",x"10",x"87"),
  1289 => (x"66",x"fc",x"c0",x"4a"),
  1290 => (x"d9",x"c8",x"c1",x"48"),
  1291 => (x"c7",x"49",x"6a",x"78"),
  1292 => (x"c0",x"51",x"74",x"81"),
  1293 => (x"c8",x"49",x"66",x"fc"),
  1294 => (x"c0",x"51",x"c1",x"81"),
  1295 => (x"c9",x"49",x"66",x"fc"),
  1296 => (x"c0",x"51",x"c0",x"81"),
  1297 => (x"ca",x"49",x"66",x"fc"),
  1298 => (x"c1",x"51",x"c0",x"81"),
  1299 => (x"6a",x"1e",x"d8",x"1e"),
  1300 => (x"e2",x"81",x"c8",x"49"),
  1301 => (x"86",x"c8",x"87",x"e1"),
  1302 => (x"48",x"66",x"c0",x"c1"),
  1303 => (x"c7",x"01",x"a8",x"c0"),
  1304 => (x"48",x"a6",x"c8",x"87"),
  1305 => (x"87",x"ce",x"78",x"c1"),
  1306 => (x"48",x"66",x"c0",x"c1"),
  1307 => (x"a6",x"d0",x"88",x"c1"),
  1308 => (x"e1",x"87",x"c3",x"58"),
  1309 => (x"a6",x"d0",x"87",x"ed"),
  1310 => (x"74",x"78",x"c2",x"48"),
  1311 => (x"cf",x"cd",x"02",x"9c"),
  1312 => (x"48",x"66",x"c8",x"87"),
  1313 => (x"a8",x"66",x"c4",x"c1"),
  1314 => (x"87",x"c4",x"cd",x"03"),
  1315 => (x"c0",x"48",x"a6",x"dc"),
  1316 => (x"c0",x"80",x"e8",x"78"),
  1317 => (x"87",x"db",x"e0",x"78"),
  1318 => (x"d0",x"c1",x"4c",x"70"),
  1319 => (x"d7",x"c2",x"05",x"ac"),
  1320 => (x"7e",x"66",x"c4",x"87"),
  1321 => (x"c8",x"87",x"ff",x"e2"),
  1322 => (x"c6",x"e0",x"58",x"a6"),
  1323 => (x"c0",x"4c",x"70",x"87"),
  1324 => (x"c1",x"05",x"ac",x"ec"),
  1325 => (x"66",x"c8",x"87",x"ed"),
  1326 => (x"c0",x"91",x"cb",x"49"),
  1327 => (x"c4",x"81",x"66",x"fc"),
  1328 => (x"4d",x"6a",x"4a",x"a1"),
  1329 => (x"c4",x"4a",x"a1",x"c8"),
  1330 => (x"c9",x"c1",x"52",x"66"),
  1331 => (x"df",x"ff",x"79",x"da"),
  1332 => (x"4c",x"70",x"87",x"e1"),
  1333 => (x"87",x"d9",x"02",x"9c"),
  1334 => (x"02",x"ac",x"fb",x"c0"),
  1335 => (x"55",x"74",x"87",x"d3"),
  1336 => (x"87",x"cf",x"df",x"ff"),
  1337 => (x"02",x"9c",x"4c",x"70"),
  1338 => (x"fb",x"c0",x"87",x"c7"),
  1339 => (x"ed",x"ff",x"05",x"ac"),
  1340 => (x"55",x"e0",x"c0",x"87"),
  1341 => (x"c0",x"55",x"c1",x"c2"),
  1342 => (x"66",x"d8",x"7d",x"97"),
  1343 => (x"05",x"a8",x"6e",x"48"),
  1344 => (x"66",x"c8",x"87",x"db"),
  1345 => (x"a8",x"66",x"cc",x"48"),
  1346 => (x"c8",x"87",x"ca",x"04"),
  1347 => (x"80",x"c1",x"48",x"66"),
  1348 => (x"c8",x"58",x"a6",x"cc"),
  1349 => (x"48",x"66",x"cc",x"87"),
  1350 => (x"a6",x"d0",x"88",x"c1"),
  1351 => (x"d2",x"de",x"ff",x"58"),
  1352 => (x"c1",x"4c",x"70",x"87"),
  1353 => (x"c8",x"05",x"ac",x"d0"),
  1354 => (x"48",x"66",x"d4",x"87"),
  1355 => (x"a6",x"d8",x"80",x"c1"),
  1356 => (x"ac",x"d0",x"c1",x"58"),
  1357 => (x"87",x"e9",x"fd",x"02"),
  1358 => (x"d8",x"48",x"66",x"c4"),
  1359 => (x"c9",x"05",x"a8",x"66"),
  1360 => (x"e0",x"c0",x"87",x"e0"),
  1361 => (x"78",x"c0",x"48",x"a6"),
  1362 => (x"fb",x"c0",x"48",x"74"),
  1363 => (x"48",x"7e",x"70",x"88"),
  1364 => (x"e2",x"c9",x"02",x"98"),
  1365 => (x"88",x"cb",x"48",x"87"),
  1366 => (x"98",x"48",x"7e",x"70"),
  1367 => (x"87",x"cd",x"c1",x"02"),
  1368 => (x"70",x"88",x"c9",x"48"),
  1369 => (x"02",x"98",x"48",x"7e"),
  1370 => (x"48",x"87",x"fe",x"c3"),
  1371 => (x"7e",x"70",x"88",x"c4"),
  1372 => (x"ce",x"02",x"98",x"48"),
  1373 => (x"88",x"c1",x"48",x"87"),
  1374 => (x"98",x"48",x"7e",x"70"),
  1375 => (x"87",x"e9",x"c3",x"02"),
  1376 => (x"dc",x"87",x"d6",x"c8"),
  1377 => (x"f0",x"c0",x"48",x"a6"),
  1378 => (x"e6",x"dc",x"ff",x"78"),
  1379 => (x"c0",x"4c",x"70",x"87"),
  1380 => (x"c0",x"02",x"ac",x"ec"),
  1381 => (x"e0",x"c0",x"87",x"c4"),
  1382 => (x"ec",x"c0",x"5c",x"a6"),
  1383 => (x"87",x"cd",x"02",x"ac"),
  1384 => (x"87",x"cf",x"dc",x"ff"),
  1385 => (x"ec",x"c0",x"4c",x"70"),
  1386 => (x"f3",x"ff",x"05",x"ac"),
  1387 => (x"ac",x"ec",x"c0",x"87"),
  1388 => (x"87",x"c4",x"c0",x"02"),
  1389 => (x"87",x"fb",x"db",x"ff"),
  1390 => (x"1e",x"ca",x"1e",x"c0"),
  1391 => (x"cb",x"49",x"66",x"d0"),
  1392 => (x"66",x"c4",x"c1",x"91"),
  1393 => (x"cc",x"80",x"71",x"48"),
  1394 => (x"66",x"c8",x"58",x"a6"),
  1395 => (x"d0",x"80",x"c4",x"48"),
  1396 => (x"66",x"cc",x"58",x"a6"),
  1397 => (x"dc",x"ff",x"49",x"bf"),
  1398 => (x"1e",x"c1",x"87",x"dd"),
  1399 => (x"66",x"d4",x"1e",x"de"),
  1400 => (x"dc",x"ff",x"49",x"bf"),
  1401 => (x"86",x"d0",x"87",x"d1"),
  1402 => (x"c0",x"48",x"49",x"70"),
  1403 => (x"e8",x"c0",x"88",x"08"),
  1404 => (x"a8",x"c0",x"58",x"a6"),
  1405 => (x"87",x"ee",x"c0",x"06"),
  1406 => (x"48",x"66",x"e4",x"c0"),
  1407 => (x"c0",x"03",x"a8",x"dd"),
  1408 => (x"66",x"c4",x"87",x"e4"),
  1409 => (x"e4",x"c0",x"49",x"bf"),
  1410 => (x"e0",x"c0",x"81",x"66"),
  1411 => (x"66",x"e4",x"c0",x"51"),
  1412 => (x"c4",x"81",x"c1",x"49"),
  1413 => (x"c2",x"81",x"bf",x"66"),
  1414 => (x"e4",x"c0",x"51",x"c1"),
  1415 => (x"81",x"c2",x"49",x"66"),
  1416 => (x"81",x"bf",x"66",x"c4"),
  1417 => (x"48",x"6e",x"51",x"c0"),
  1418 => (x"78",x"d9",x"c8",x"c1"),
  1419 => (x"81",x"c8",x"49",x"6e"),
  1420 => (x"6e",x"51",x"66",x"d0"),
  1421 => (x"d4",x"81",x"c9",x"49"),
  1422 => (x"49",x"6e",x"51",x"66"),
  1423 => (x"66",x"dc",x"81",x"ca"),
  1424 => (x"48",x"66",x"d0",x"51"),
  1425 => (x"a6",x"d4",x"80",x"c1"),
  1426 => (x"48",x"66",x"c8",x"58"),
  1427 => (x"04",x"a8",x"66",x"cc"),
  1428 => (x"c8",x"87",x"cb",x"c0"),
  1429 => (x"80",x"c1",x"48",x"66"),
  1430 => (x"c5",x"58",x"a6",x"cc"),
  1431 => (x"66",x"cc",x"87",x"d9"),
  1432 => (x"d0",x"88",x"c1",x"48"),
  1433 => (x"ce",x"c5",x"58",x"a6"),
  1434 => (x"f9",x"db",x"ff",x"87"),
  1435 => (x"a6",x"e8",x"c0",x"87"),
  1436 => (x"f1",x"db",x"ff",x"58"),
  1437 => (x"a6",x"e0",x"c0",x"87"),
  1438 => (x"a8",x"ec",x"c0",x"58"),
  1439 => (x"87",x"ca",x"c0",x"05"),
  1440 => (x"c0",x"48",x"a6",x"dc"),
  1441 => (x"c0",x"78",x"66",x"e4"),
  1442 => (x"d8",x"ff",x"87",x"c4"),
  1443 => (x"66",x"c8",x"87",x"e5"),
  1444 => (x"c0",x"91",x"cb",x"49"),
  1445 => (x"71",x"48",x"66",x"fc"),
  1446 => (x"4a",x"7e",x"70",x"80"),
  1447 => (x"49",x"6e",x"82",x"c8"),
  1448 => (x"e4",x"c0",x"81",x"ca"),
  1449 => (x"66",x"dc",x"51",x"66"),
  1450 => (x"c0",x"81",x"c1",x"49"),
  1451 => (x"c1",x"89",x"66",x"e4"),
  1452 => (x"70",x"30",x"71",x"48"),
  1453 => (x"71",x"89",x"c1",x"49"),
  1454 => (x"ed",x"c2",x"7a",x"97"),
  1455 => (x"c0",x"49",x"bf",x"f8"),
  1456 => (x"97",x"29",x"66",x"e4"),
  1457 => (x"71",x"48",x"4a",x"6a"),
  1458 => (x"a6",x"ec",x"c0",x"98"),
  1459 => (x"c4",x"49",x"6e",x"58"),
  1460 => (x"d8",x"4d",x"69",x"81"),
  1461 => (x"66",x"c4",x"48",x"66"),
  1462 => (x"c8",x"c0",x"02",x"a8"),
  1463 => (x"48",x"a6",x"c4",x"87"),
  1464 => (x"c5",x"c0",x"78",x"c0"),
  1465 => (x"48",x"a6",x"c4",x"87"),
  1466 => (x"66",x"c4",x"78",x"c1"),
  1467 => (x"1e",x"e0",x"c0",x"1e"),
  1468 => (x"d8",x"ff",x"49",x"75"),
  1469 => (x"86",x"c8",x"87",x"c1"),
  1470 => (x"b7",x"c0",x"4c",x"70"),
  1471 => (x"d4",x"c1",x"06",x"ac"),
  1472 => (x"c0",x"85",x"74",x"87"),
  1473 => (x"89",x"74",x"49",x"e0"),
  1474 => (x"e0",x"c1",x"4b",x"75"),
  1475 => (x"fe",x"71",x"4a",x"d2"),
  1476 => (x"c2",x"87",x"d4",x"e6"),
  1477 => (x"66",x"e0",x"c0",x"85"),
  1478 => (x"c0",x"80",x"c1",x"48"),
  1479 => (x"c0",x"58",x"a6",x"e4"),
  1480 => (x"c1",x"49",x"66",x"e8"),
  1481 => (x"02",x"a9",x"70",x"81"),
  1482 => (x"c4",x"87",x"c8",x"c0"),
  1483 => (x"78",x"c0",x"48",x"a6"),
  1484 => (x"c4",x"87",x"c5",x"c0"),
  1485 => (x"78",x"c1",x"48",x"a6"),
  1486 => (x"c2",x"1e",x"66",x"c4"),
  1487 => (x"e0",x"c0",x"49",x"a4"),
  1488 => (x"70",x"88",x"71",x"48"),
  1489 => (x"49",x"75",x"1e",x"49"),
  1490 => (x"87",x"eb",x"d6",x"ff"),
  1491 => (x"b7",x"c0",x"86",x"c8"),
  1492 => (x"c0",x"ff",x"01",x"a8"),
  1493 => (x"66",x"e0",x"c0",x"87"),
  1494 => (x"87",x"d1",x"c0",x"02"),
  1495 => (x"81",x"c9",x"49",x"6e"),
  1496 => (x"51",x"66",x"e0",x"c0"),
  1497 => (x"ca",x"c1",x"48",x"6e"),
  1498 => (x"cc",x"c0",x"78",x"ea"),
  1499 => (x"c9",x"49",x"6e",x"87"),
  1500 => (x"6e",x"51",x"c2",x"81"),
  1501 => (x"d6",x"cc",x"c1",x"48"),
  1502 => (x"48",x"66",x"c8",x"78"),
  1503 => (x"04",x"a8",x"66",x"cc"),
  1504 => (x"c8",x"87",x"cb",x"c0"),
  1505 => (x"80",x"c1",x"48",x"66"),
  1506 => (x"c0",x"58",x"a6",x"cc"),
  1507 => (x"66",x"cc",x"87",x"e9"),
  1508 => (x"d0",x"88",x"c1",x"48"),
  1509 => (x"de",x"c0",x"58",x"a6"),
  1510 => (x"c6",x"d5",x"ff",x"87"),
  1511 => (x"c0",x"4c",x"70",x"87"),
  1512 => (x"c6",x"c1",x"87",x"d5"),
  1513 => (x"c8",x"c0",x"05",x"ac"),
  1514 => (x"48",x"66",x"d0",x"87"),
  1515 => (x"a6",x"d4",x"80",x"c1"),
  1516 => (x"ee",x"d4",x"ff",x"58"),
  1517 => (x"d4",x"4c",x"70",x"87"),
  1518 => (x"80",x"c1",x"48",x"66"),
  1519 => (x"74",x"58",x"a6",x"d8"),
  1520 => (x"cb",x"c0",x"02",x"9c"),
  1521 => (x"48",x"66",x"c8",x"87"),
  1522 => (x"a8",x"66",x"c4",x"c1"),
  1523 => (x"87",x"fc",x"f2",x"04"),
  1524 => (x"87",x"c6",x"d4",x"ff"),
  1525 => (x"c7",x"48",x"66",x"c8"),
  1526 => (x"e5",x"c0",x"03",x"a8"),
  1527 => (x"cc",x"ea",x"c2",x"87"),
  1528 => (x"c8",x"78",x"c0",x"48"),
  1529 => (x"91",x"cb",x"49",x"66"),
  1530 => (x"81",x"66",x"fc",x"c0"),
  1531 => (x"6a",x"4a",x"a1",x"c4"),
  1532 => (x"79",x"52",x"c0",x"4a"),
  1533 => (x"c1",x"48",x"66",x"c8"),
  1534 => (x"58",x"a6",x"cc",x"80"),
  1535 => (x"ff",x"04",x"a8",x"c7"),
  1536 => (x"d4",x"ff",x"87",x"db"),
  1537 => (x"d6",x"de",x"ff",x"8e"),
  1538 => (x"61",x"6f",x"4c",x"87"),
  1539 => (x"2e",x"2a",x"20",x"64"),
  1540 => (x"20",x"3a",x"00",x"20"),
  1541 => (x"1e",x"73",x"1e",x"00"),
  1542 => (x"02",x"9b",x"4b",x"71"),
  1543 => (x"ea",x"c2",x"87",x"c6"),
  1544 => (x"78",x"c0",x"48",x"c8"),
  1545 => (x"ea",x"c2",x"1e",x"c7"),
  1546 => (x"c1",x"1e",x"bf",x"c8"),
  1547 => (x"c2",x"1e",x"f0",x"e3"),
  1548 => (x"49",x"bf",x"f0",x"e9"),
  1549 => (x"cc",x"87",x"ff",x"ed"),
  1550 => (x"f0",x"e9",x"c2",x"86"),
  1551 => (x"c1",x"e9",x"49",x"bf"),
  1552 => (x"02",x"9b",x"73",x"87"),
  1553 => (x"e3",x"c1",x"87",x"c8"),
  1554 => (x"e2",x"c0",x"49",x"f0"),
  1555 => (x"dd",x"ff",x"87",x"da"),
  1556 => (x"c7",x"1e",x"87",x"d1"),
  1557 => (x"49",x"c1",x"87",x"d1"),
  1558 => (x"fe",x"87",x"fa",x"fe"),
  1559 => (x"70",x"87",x"f8",x"e9"),
  1560 => (x"87",x"cd",x"02",x"98"),
  1561 => (x"87",x"f2",x"f2",x"fe"),
  1562 => (x"c4",x"02",x"98",x"70"),
  1563 => (x"c2",x"4a",x"c1",x"87"),
  1564 => (x"72",x"4a",x"c0",x"87"),
  1565 => (x"87",x"ce",x"05",x"9a"),
  1566 => (x"e2",x"c1",x"1e",x"c0"),
  1567 => (x"ef",x"c0",x"49",x"e3"),
  1568 => (x"86",x"c4",x"87",x"d2"),
  1569 => (x"1e",x"c0",x"87",x"fe"),
  1570 => (x"49",x"ee",x"e2",x"c1"),
  1571 => (x"87",x"c4",x"ef",x"c0"),
  1572 => (x"f8",x"c0",x"1e",x"c0"),
  1573 => (x"49",x"70",x"87",x"e1"),
  1574 => (x"87",x"f8",x"ee",x"c0"),
  1575 => (x"f8",x"87",x"c7",x"c3"),
  1576 => (x"53",x"4f",x"26",x"8e"),
  1577 => (x"61",x"66",x"20",x"44"),
  1578 => (x"64",x"65",x"6c",x"69"),
  1579 => (x"6f",x"42",x"00",x"2e"),
  1580 => (x"6e",x"69",x"74",x"6f"),
  1581 => (x"2e",x"2e",x"2e",x"67"),
  1582 => (x"e5",x"c0",x"1e",x"00"),
  1583 => (x"f2",x"c0",x"87",x"e7"),
  1584 => (x"87",x"f6",x"87",x"dd"),
  1585 => (x"c2",x"1e",x"4f",x"26"),
  1586 => (x"c0",x"48",x"c8",x"ea"),
  1587 => (x"f0",x"e9",x"c2",x"78"),
  1588 => (x"fd",x"78",x"c0",x"48"),
  1589 => (x"87",x"e1",x"87",x"fc"),
  1590 => (x"4f",x"26",x"48",x"c0"),
  1591 => (x"00",x"01",x"00",x"00"),
  1592 => (x"20",x"80",x"00",x"00"),
  1593 => (x"74",x"69",x"78",x"45"),
  1594 => (x"42",x"20",x"80",x"00"),
  1595 => (x"00",x"6b",x"63",x"61"),
  1596 => (x"00",x"00",x"10",x"26"),
  1597 => (x"00",x"00",x"2a",x"9c"),
  1598 => (x"26",x"00",x"00",x"00"),
  1599 => (x"ba",x"00",x"00",x"10"),
  1600 => (x"00",x"00",x"00",x"2a"),
  1601 => (x"10",x"26",x"00",x"00"),
  1602 => (x"2a",x"d8",x"00",x"00"),
  1603 => (x"00",x"00",x"00",x"00"),
  1604 => (x"00",x"10",x"26",x"00"),
  1605 => (x"00",x"2a",x"f6",x"00"),
  1606 => (x"00",x"00",x"00",x"00"),
  1607 => (x"00",x"00",x"10",x"26"),
  1608 => (x"00",x"00",x"2b",x"14"),
  1609 => (x"26",x"00",x"00",x"00"),
  1610 => (x"32",x"00",x"00",x"10"),
  1611 => (x"00",x"00",x"00",x"2b"),
  1612 => (x"10",x"26",x"00",x"00"),
  1613 => (x"2b",x"50",x"00",x"00"),
  1614 => (x"00",x"00",x"00",x"00"),
  1615 => (x"00",x"12",x"5a",x"00"),
  1616 => (x"00",x"00",x"00",x"00"),
  1617 => (x"00",x"00",x"00",x"00"),
  1618 => (x"00",x"00",x"13",x"27"),
  1619 => (x"00",x"00",x"00",x"00"),
  1620 => (x"1e",x"00",x"00",x"00"),
  1621 => (x"c0",x"48",x"f0",x"fe"),
  1622 => (x"79",x"09",x"cd",x"78"),
  1623 => (x"1e",x"4f",x"26",x"09"),
  1624 => (x"48",x"bf",x"f0",x"fe"),
  1625 => (x"fe",x"1e",x"4f",x"26"),
  1626 => (x"78",x"c1",x"48",x"f0"),
  1627 => (x"fe",x"1e",x"4f",x"26"),
  1628 => (x"78",x"c0",x"48",x"f0"),
  1629 => (x"71",x"1e",x"4f",x"26"),
  1630 => (x"51",x"52",x"c0",x"4a"),
  1631 => (x"5e",x"0e",x"4f",x"26"),
  1632 => (x"0e",x"5d",x"5c",x"5b"),
  1633 => (x"4d",x"71",x"86",x"f4"),
  1634 => (x"c1",x"7e",x"6d",x"97"),
  1635 => (x"6c",x"97",x"4c",x"a5"),
  1636 => (x"58",x"a6",x"c8",x"48"),
  1637 => (x"66",x"c4",x"48",x"6e"),
  1638 => (x"87",x"c5",x"05",x"a8"),
  1639 => (x"e6",x"c0",x"48",x"ff"),
  1640 => (x"87",x"ca",x"ff",x"87"),
  1641 => (x"97",x"49",x"a5",x"c2"),
  1642 => (x"a3",x"71",x"4b",x"6c"),
  1643 => (x"4b",x"6b",x"97",x"4b"),
  1644 => (x"6e",x"7e",x"6c",x"97"),
  1645 => (x"c8",x"80",x"c1",x"48"),
  1646 => (x"98",x"c7",x"58",x"a6"),
  1647 => (x"70",x"58",x"a6",x"cc"),
  1648 => (x"e1",x"fe",x"7c",x"97"),
  1649 => (x"f4",x"48",x"73",x"87"),
  1650 => (x"26",x"4d",x"26",x"8e"),
  1651 => (x"26",x"4b",x"26",x"4c"),
  1652 => (x"5b",x"5e",x"0e",x"4f"),
  1653 => (x"86",x"f4",x"0e",x"5c"),
  1654 => (x"66",x"d8",x"4c",x"71"),
  1655 => (x"9a",x"ff",x"c3",x"4a"),
  1656 => (x"97",x"4b",x"a4",x"c2"),
  1657 => (x"a1",x"73",x"49",x"6c"),
  1658 => (x"97",x"51",x"72",x"49"),
  1659 => (x"48",x"6e",x"7e",x"6c"),
  1660 => (x"a6",x"c8",x"80",x"c1"),
  1661 => (x"cc",x"98",x"c7",x"58"),
  1662 => (x"54",x"70",x"58",x"a6"),
  1663 => (x"ca",x"ff",x"8e",x"f4"),
  1664 => (x"fd",x"1e",x"1e",x"87"),
  1665 => (x"bf",x"e0",x"87",x"e8"),
  1666 => (x"e0",x"c0",x"49",x"4a"),
  1667 => (x"cb",x"02",x"99",x"c0"),
  1668 => (x"c2",x"1e",x"72",x"87"),
  1669 => (x"fe",x"49",x"ee",x"ed"),
  1670 => (x"86",x"c4",x"87",x"f7"),
  1671 => (x"70",x"87",x"c0",x"fd"),
  1672 => (x"87",x"c2",x"fd",x"7e"),
  1673 => (x"1e",x"4f",x"26",x"26"),
  1674 => (x"49",x"ee",x"ed",x"c2"),
  1675 => (x"c1",x"87",x"c7",x"fd"),
  1676 => (x"fc",x"49",x"c1",x"e8"),
  1677 => (x"f7",x"c3",x"87",x"dd"),
  1678 => (x"0e",x"4f",x"26",x"87"),
  1679 => (x"5d",x"5c",x"5b",x"5e"),
  1680 => (x"c2",x"4d",x"71",x"0e"),
  1681 => (x"fc",x"49",x"ee",x"ed"),
  1682 => (x"4b",x"70",x"87",x"f4"),
  1683 => (x"04",x"ab",x"b7",x"c0"),
  1684 => (x"c3",x"87",x"c2",x"c3"),
  1685 => (x"c9",x"05",x"ab",x"f0"),
  1686 => (x"df",x"ec",x"c1",x"87"),
  1687 => (x"c2",x"78",x"c1",x"48"),
  1688 => (x"e0",x"c3",x"87",x"e3"),
  1689 => (x"87",x"c9",x"05",x"ab"),
  1690 => (x"48",x"e3",x"ec",x"c1"),
  1691 => (x"d4",x"c2",x"78",x"c1"),
  1692 => (x"e3",x"ec",x"c1",x"87"),
  1693 => (x"87",x"c6",x"02",x"bf"),
  1694 => (x"4c",x"a3",x"c0",x"c2"),
  1695 => (x"4c",x"73",x"87",x"c2"),
  1696 => (x"bf",x"df",x"ec",x"c1"),
  1697 => (x"87",x"e0",x"c0",x"02"),
  1698 => (x"b7",x"c4",x"49",x"74"),
  1699 => (x"ed",x"c1",x"91",x"29"),
  1700 => (x"4a",x"74",x"81",x"ff"),
  1701 => (x"92",x"c2",x"9a",x"cf"),
  1702 => (x"30",x"72",x"48",x"c1"),
  1703 => (x"ba",x"ff",x"4a",x"70"),
  1704 => (x"98",x"69",x"48",x"72"),
  1705 => (x"87",x"db",x"79",x"70"),
  1706 => (x"b7",x"c4",x"49",x"74"),
  1707 => (x"ed",x"c1",x"91",x"29"),
  1708 => (x"4a",x"74",x"81",x"ff"),
  1709 => (x"92",x"c2",x"9a",x"cf"),
  1710 => (x"30",x"72",x"48",x"c3"),
  1711 => (x"69",x"48",x"4a",x"70"),
  1712 => (x"75",x"79",x"70",x"b0"),
  1713 => (x"f0",x"c0",x"05",x"9d"),
  1714 => (x"48",x"d0",x"ff",x"87"),
  1715 => (x"ff",x"78",x"e1",x"c8"),
  1716 => (x"78",x"c5",x"48",x"d4"),
  1717 => (x"bf",x"e3",x"ec",x"c1"),
  1718 => (x"c3",x"87",x"c3",x"02"),
  1719 => (x"ec",x"c1",x"78",x"e0"),
  1720 => (x"c6",x"02",x"bf",x"df"),
  1721 => (x"48",x"d4",x"ff",x"87"),
  1722 => (x"ff",x"78",x"f0",x"c3"),
  1723 => (x"0b",x"7b",x"0b",x"d4"),
  1724 => (x"c8",x"48",x"d0",x"ff"),
  1725 => (x"e0",x"c0",x"78",x"e1"),
  1726 => (x"e3",x"ec",x"c1",x"78"),
  1727 => (x"c1",x"78",x"c0",x"48"),
  1728 => (x"c0",x"48",x"df",x"ec"),
  1729 => (x"ee",x"ed",x"c2",x"78"),
  1730 => (x"87",x"f2",x"f9",x"49"),
  1731 => (x"b7",x"c0",x"4b",x"70"),
  1732 => (x"fe",x"fc",x"03",x"ab"),
  1733 => (x"26",x"48",x"c0",x"87"),
  1734 => (x"26",x"4c",x"26",x"4d"),
  1735 => (x"00",x"4f",x"26",x"4b"),
  1736 => (x"00",x"00",x"00",x"00"),
  1737 => (x"1e",x"00",x"00",x"00"),
  1738 => (x"fc",x"49",x"4a",x"71"),
  1739 => (x"4f",x"26",x"87",x"cd"),
  1740 => (x"72",x"4a",x"c0",x"1e"),
  1741 => (x"c1",x"91",x"c4",x"49"),
  1742 => (x"c0",x"81",x"ff",x"ed"),
  1743 => (x"d0",x"82",x"c1",x"79"),
  1744 => (x"ee",x"04",x"aa",x"b7"),
  1745 => (x"0e",x"4f",x"26",x"87"),
  1746 => (x"5d",x"5c",x"5b",x"5e"),
  1747 => (x"f8",x"4d",x"71",x"0e"),
  1748 => (x"4a",x"75",x"87",x"dc"),
  1749 => (x"92",x"2a",x"b7",x"c4"),
  1750 => (x"82",x"ff",x"ed",x"c1"),
  1751 => (x"9c",x"cf",x"4c",x"75"),
  1752 => (x"49",x"6a",x"94",x"c2"),
  1753 => (x"c3",x"2b",x"74",x"4b"),
  1754 => (x"74",x"48",x"c2",x"9b"),
  1755 => (x"ff",x"4c",x"70",x"30"),
  1756 => (x"71",x"48",x"74",x"bc"),
  1757 => (x"f7",x"7a",x"70",x"98"),
  1758 => (x"48",x"73",x"87",x"ec"),
  1759 => (x"00",x"87",x"d8",x"fe"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"00",x"00"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"1e",x"00",x"00",x"00"),
  1776 => (x"c8",x"48",x"d0",x"ff"),
  1777 => (x"48",x"71",x"78",x"e1"),
  1778 => (x"78",x"08",x"d4",x"ff"),
  1779 => (x"ff",x"1e",x"4f",x"26"),
  1780 => (x"e1",x"c8",x"48",x"d0"),
  1781 => (x"ff",x"48",x"71",x"78"),
  1782 => (x"c4",x"78",x"08",x"d4"),
  1783 => (x"d4",x"ff",x"48",x"66"),
  1784 => (x"4f",x"26",x"78",x"08"),
  1785 => (x"c4",x"4a",x"71",x"1e"),
  1786 => (x"72",x"1e",x"49",x"66"),
  1787 => (x"87",x"de",x"ff",x"49"),
  1788 => (x"c0",x"48",x"d0",x"ff"),
  1789 => (x"26",x"26",x"78",x"e0"),
  1790 => (x"1e",x"73",x"1e",x"4f"),
  1791 => (x"66",x"c8",x"4b",x"71"),
  1792 => (x"4a",x"73",x"1e",x"49"),
  1793 => (x"49",x"a2",x"e0",x"c1"),
  1794 => (x"26",x"87",x"d9",x"ff"),
  1795 => (x"4d",x"26",x"87",x"c4"),
  1796 => (x"4b",x"26",x"4c",x"26"),
  1797 => (x"ff",x"1e",x"4f",x"26"),
  1798 => (x"ff",x"c3",x"4a",x"d4"),
  1799 => (x"48",x"d0",x"ff",x"7a"),
  1800 => (x"de",x"78",x"e1",x"c0"),
  1801 => (x"f8",x"ed",x"c2",x"7a"),
  1802 => (x"48",x"49",x"7a",x"bf"),
  1803 => (x"7a",x"70",x"28",x"c8"),
  1804 => (x"28",x"d0",x"48",x"71"),
  1805 => (x"48",x"71",x"7a",x"70"),
  1806 => (x"7a",x"70",x"28",x"d8"),
  1807 => (x"c0",x"48",x"d0",x"ff"),
  1808 => (x"4f",x"26",x"78",x"e0"),
  1809 => (x"48",x"d0",x"ff",x"1e"),
  1810 => (x"71",x"78",x"c9",x"c8"),
  1811 => (x"08",x"d4",x"ff",x"48"),
  1812 => (x"1e",x"4f",x"26",x"78"),
  1813 => (x"eb",x"49",x"4a",x"71"),
  1814 => (x"48",x"d0",x"ff",x"87"),
  1815 => (x"4f",x"26",x"78",x"c8"),
  1816 => (x"71",x"1e",x"73",x"1e"),
  1817 => (x"c8",x"ee",x"c2",x"4b"),
  1818 => (x"87",x"c3",x"02",x"bf"),
  1819 => (x"ff",x"87",x"eb",x"c2"),
  1820 => (x"c9",x"c8",x"48",x"d0"),
  1821 => (x"c0",x"48",x"73",x"78"),
  1822 => (x"d4",x"ff",x"b0",x"e0"),
  1823 => (x"ed",x"c2",x"78",x"08"),
  1824 => (x"78",x"c0",x"48",x"fc"),
  1825 => (x"c5",x"02",x"66",x"c8"),
  1826 => (x"49",x"ff",x"c3",x"87"),
  1827 => (x"49",x"c0",x"87",x"c2"),
  1828 => (x"59",x"c4",x"ee",x"c2"),
  1829 => (x"c6",x"02",x"66",x"cc"),
  1830 => (x"d5",x"d5",x"c5",x"87"),
  1831 => (x"cf",x"87",x"c4",x"4a"),
  1832 => (x"c2",x"4a",x"ff",x"ff"),
  1833 => (x"c2",x"5a",x"c8",x"ee"),
  1834 => (x"c1",x"48",x"c8",x"ee"),
  1835 => (x"26",x"87",x"c4",x"78"),
  1836 => (x"26",x"4c",x"26",x"4d"),
  1837 => (x"0e",x"4f",x"26",x"4b"),
  1838 => (x"5d",x"5c",x"5b",x"5e"),
  1839 => (x"c2",x"4a",x"71",x"0e"),
  1840 => (x"4c",x"bf",x"c4",x"ee"),
  1841 => (x"cb",x"02",x"9a",x"72"),
  1842 => (x"91",x"c8",x"49",x"87"),
  1843 => (x"4b",x"d6",x"f1",x"c1"),
  1844 => (x"87",x"c4",x"83",x"71"),
  1845 => (x"4b",x"d6",x"f5",x"c1"),
  1846 => (x"49",x"13",x"4d",x"c0"),
  1847 => (x"ee",x"c2",x"99",x"74"),
  1848 => (x"71",x"48",x"bf",x"c0"),
  1849 => (x"08",x"d4",x"ff",x"b8"),
  1850 => (x"2c",x"b7",x"c1",x"78"),
  1851 => (x"ad",x"b7",x"c8",x"85"),
  1852 => (x"c2",x"87",x"e7",x"04"),
  1853 => (x"48",x"bf",x"fc",x"ed"),
  1854 => (x"ee",x"c2",x"80",x"c8"),
  1855 => (x"ee",x"fe",x"58",x"c0"),
  1856 => (x"1e",x"73",x"1e",x"87"),
  1857 => (x"4a",x"13",x"4b",x"71"),
  1858 => (x"87",x"cb",x"02",x"9a"),
  1859 => (x"e6",x"fe",x"49",x"72"),
  1860 => (x"9a",x"4a",x"13",x"87"),
  1861 => (x"fe",x"87",x"f5",x"05"),
  1862 => (x"c2",x"1e",x"87",x"d9"),
  1863 => (x"49",x"bf",x"fc",x"ed"),
  1864 => (x"48",x"fc",x"ed",x"c2"),
  1865 => (x"c4",x"78",x"a1",x"c1"),
  1866 => (x"03",x"a9",x"b7",x"c0"),
  1867 => (x"d4",x"ff",x"87",x"db"),
  1868 => (x"c0",x"ee",x"c2",x"48"),
  1869 => (x"ed",x"c2",x"78",x"bf"),
  1870 => (x"c2",x"49",x"bf",x"fc"),
  1871 => (x"c1",x"48",x"fc",x"ed"),
  1872 => (x"c0",x"c4",x"78",x"a1"),
  1873 => (x"e5",x"04",x"a9",x"b7"),
  1874 => (x"48",x"d0",x"ff",x"87"),
  1875 => (x"ee",x"c2",x"78",x"c8"),
  1876 => (x"78",x"c0",x"48",x"c8"),
  1877 => (x"00",x"00",x"4f",x"26"),
  1878 => (x"00",x"00",x"00",x"00"),
  1879 => (x"00",x"00",x"00",x"00"),
  1880 => (x"00",x"5f",x"5f",x"00"),
  1881 => (x"03",x"00",x"00",x"00"),
  1882 => (x"03",x"03",x"00",x"03"),
  1883 => (x"7f",x"14",x"00",x"00"),
  1884 => (x"7f",x"7f",x"14",x"7f"),
  1885 => (x"24",x"00",x"00",x"14"),
  1886 => (x"3a",x"6b",x"6b",x"2e"),
  1887 => (x"6a",x"4c",x"00",x"12"),
  1888 => (x"56",x"6c",x"18",x"36"),
  1889 => (x"7e",x"30",x"00",x"32"),
  1890 => (x"3a",x"77",x"59",x"4f"),
  1891 => (x"00",x"00",x"40",x"68"),
  1892 => (x"00",x"03",x"07",x"04"),
  1893 => (x"00",x"00",x"00",x"00"),
  1894 => (x"41",x"63",x"3e",x"1c"),
  1895 => (x"00",x"00",x"00",x"00"),
  1896 => (x"1c",x"3e",x"63",x"41"),
  1897 => (x"2a",x"08",x"00",x"00"),
  1898 => (x"3e",x"1c",x"1c",x"3e"),
  1899 => (x"08",x"00",x"08",x"2a"),
  1900 => (x"08",x"3e",x"3e",x"08"),
  1901 => (x"00",x"00",x"00",x"08"),
  1902 => (x"00",x"60",x"e0",x"80"),
  1903 => (x"08",x"00",x"00",x"00"),
  1904 => (x"08",x"08",x"08",x"08"),
  1905 => (x"00",x"00",x"00",x"08"),
  1906 => (x"00",x"60",x"60",x"00"),
  1907 => (x"60",x"40",x"00",x"00"),
  1908 => (x"06",x"0c",x"18",x"30"),
  1909 => (x"3e",x"00",x"01",x"03"),
  1910 => (x"7f",x"4d",x"59",x"7f"),
  1911 => (x"04",x"00",x"00",x"3e"),
  1912 => (x"00",x"7f",x"7f",x"06"),
  1913 => (x"42",x"00",x"00",x"00"),
  1914 => (x"4f",x"59",x"71",x"63"),
  1915 => (x"22",x"00",x"00",x"46"),
  1916 => (x"7f",x"49",x"49",x"63"),
  1917 => (x"1c",x"18",x"00",x"36"),
  1918 => (x"7f",x"7f",x"13",x"16"),
  1919 => (x"27",x"00",x"00",x"10"),
  1920 => (x"7d",x"45",x"45",x"67"),
  1921 => (x"3c",x"00",x"00",x"39"),
  1922 => (x"79",x"49",x"4b",x"7e"),
  1923 => (x"01",x"00",x"00",x"30"),
  1924 => (x"0f",x"79",x"71",x"01"),
  1925 => (x"36",x"00",x"00",x"07"),
  1926 => (x"7f",x"49",x"49",x"7f"),
  1927 => (x"06",x"00",x"00",x"36"),
  1928 => (x"3f",x"69",x"49",x"4f"),
  1929 => (x"00",x"00",x"00",x"1e"),
  1930 => (x"00",x"66",x"66",x"00"),
  1931 => (x"00",x"00",x"00",x"00"),
  1932 => (x"00",x"66",x"e6",x"80"),
  1933 => (x"08",x"00",x"00",x"00"),
  1934 => (x"22",x"14",x"14",x"08"),
  1935 => (x"14",x"00",x"00",x"22"),
  1936 => (x"14",x"14",x"14",x"14"),
  1937 => (x"22",x"00",x"00",x"14"),
  1938 => (x"08",x"14",x"14",x"22"),
  1939 => (x"02",x"00",x"00",x"08"),
  1940 => (x"0f",x"59",x"51",x"03"),
  1941 => (x"7f",x"3e",x"00",x"06"),
  1942 => (x"1f",x"55",x"5d",x"41"),
  1943 => (x"7e",x"00",x"00",x"1e"),
  1944 => (x"7f",x"09",x"09",x"7f"),
  1945 => (x"7f",x"00",x"00",x"7e"),
  1946 => (x"7f",x"49",x"49",x"7f"),
  1947 => (x"1c",x"00",x"00",x"36"),
  1948 => (x"41",x"41",x"63",x"3e"),
  1949 => (x"7f",x"00",x"00",x"41"),
  1950 => (x"3e",x"63",x"41",x"7f"),
  1951 => (x"7f",x"00",x"00",x"1c"),
  1952 => (x"41",x"49",x"49",x"7f"),
  1953 => (x"7f",x"00",x"00",x"41"),
  1954 => (x"01",x"09",x"09",x"7f"),
  1955 => (x"3e",x"00",x"00",x"01"),
  1956 => (x"7b",x"49",x"41",x"7f"),
  1957 => (x"7f",x"00",x"00",x"7a"),
  1958 => (x"7f",x"08",x"08",x"7f"),
  1959 => (x"00",x"00",x"00",x"7f"),
  1960 => (x"41",x"7f",x"7f",x"41"),
  1961 => (x"20",x"00",x"00",x"00"),
  1962 => (x"7f",x"40",x"40",x"60"),
  1963 => (x"7f",x"7f",x"00",x"3f"),
  1964 => (x"63",x"36",x"1c",x"08"),
  1965 => (x"7f",x"00",x"00",x"41"),
  1966 => (x"40",x"40",x"40",x"7f"),
  1967 => (x"7f",x"7f",x"00",x"40"),
  1968 => (x"7f",x"06",x"0c",x"06"),
  1969 => (x"7f",x"7f",x"00",x"7f"),
  1970 => (x"7f",x"18",x"0c",x"06"),
  1971 => (x"3e",x"00",x"00",x"7f"),
  1972 => (x"7f",x"41",x"41",x"7f"),
  1973 => (x"7f",x"00",x"00",x"3e"),
  1974 => (x"0f",x"09",x"09",x"7f"),
  1975 => (x"7f",x"3e",x"00",x"06"),
  1976 => (x"7e",x"7f",x"61",x"41"),
  1977 => (x"7f",x"00",x"00",x"40"),
  1978 => (x"7f",x"19",x"09",x"7f"),
  1979 => (x"26",x"00",x"00",x"66"),
  1980 => (x"7b",x"59",x"4d",x"6f"),
  1981 => (x"01",x"00",x"00",x"32"),
  1982 => (x"01",x"7f",x"7f",x"01"),
  1983 => (x"3f",x"00",x"00",x"01"),
  1984 => (x"7f",x"40",x"40",x"7f"),
  1985 => (x"0f",x"00",x"00",x"3f"),
  1986 => (x"3f",x"70",x"70",x"3f"),
  1987 => (x"7f",x"7f",x"00",x"0f"),
  1988 => (x"7f",x"30",x"18",x"30"),
  1989 => (x"63",x"41",x"00",x"7f"),
  1990 => (x"36",x"1c",x"1c",x"36"),
  1991 => (x"03",x"01",x"41",x"63"),
  1992 => (x"06",x"7c",x"7c",x"06"),
  1993 => (x"71",x"61",x"01",x"03"),
  1994 => (x"43",x"47",x"4d",x"59"),
  1995 => (x"00",x"00",x"00",x"41"),
  1996 => (x"41",x"41",x"7f",x"7f"),
  1997 => (x"03",x"01",x"00",x"00"),
  1998 => (x"30",x"18",x"0c",x"06"),
  1999 => (x"00",x"00",x"40",x"60"),
  2000 => (x"7f",x"7f",x"41",x"41"),
  2001 => (x"0c",x"08",x"00",x"00"),
  2002 => (x"0c",x"06",x"03",x"06"),
  2003 => (x"80",x"80",x"00",x"08"),
  2004 => (x"80",x"80",x"80",x"80"),
  2005 => (x"00",x"00",x"00",x"80"),
  2006 => (x"04",x"07",x"03",x"00"),
  2007 => (x"20",x"00",x"00",x"00"),
  2008 => (x"7c",x"54",x"54",x"74"),
  2009 => (x"7f",x"00",x"00",x"78"),
  2010 => (x"7c",x"44",x"44",x"7f"),
  2011 => (x"38",x"00",x"00",x"38"),
  2012 => (x"44",x"44",x"44",x"7c"),
  2013 => (x"38",x"00",x"00",x"00"),
  2014 => (x"7f",x"44",x"44",x"7c"),
  2015 => (x"38",x"00",x"00",x"7f"),
  2016 => (x"5c",x"54",x"54",x"7c"),
  2017 => (x"04",x"00",x"00",x"18"),
  2018 => (x"05",x"05",x"7f",x"7e"),
  2019 => (x"18",x"00",x"00",x"00"),
  2020 => (x"fc",x"a4",x"a4",x"bc"),
  2021 => (x"7f",x"00",x"00",x"7c"),
  2022 => (x"7c",x"04",x"04",x"7f"),
  2023 => (x"00",x"00",x"00",x"78"),
  2024 => (x"40",x"7d",x"3d",x"00"),
  2025 => (x"80",x"00",x"00",x"00"),
  2026 => (x"7d",x"fd",x"80",x"80"),
  2027 => (x"7f",x"00",x"00",x"00"),
  2028 => (x"6c",x"38",x"10",x"7f"),
  2029 => (x"00",x"00",x"00",x"44"),
  2030 => (x"40",x"7f",x"3f",x"00"),
  2031 => (x"7c",x"7c",x"00",x"00"),
  2032 => (x"7c",x"0c",x"18",x"0c"),
  2033 => (x"7c",x"00",x"00",x"78"),
  2034 => (x"7c",x"04",x"04",x"7c"),
  2035 => (x"38",x"00",x"00",x"78"),
  2036 => (x"7c",x"44",x"44",x"7c"),
  2037 => (x"fc",x"00",x"00",x"38"),
  2038 => (x"3c",x"24",x"24",x"fc"),
  2039 => (x"18",x"00",x"00",x"18"),
  2040 => (x"fc",x"24",x"24",x"3c"),
  2041 => (x"7c",x"00",x"00",x"fc"),
  2042 => (x"0c",x"04",x"04",x"7c"),
  2043 => (x"48",x"00",x"00",x"08"),
  2044 => (x"74",x"54",x"54",x"5c"),
  2045 => (x"04",x"00",x"00",x"20"),
  2046 => (x"44",x"44",x"7f",x"3f"),
  2047 => (x"3c",x"00",x"00",x"00"),
  2048 => (x"7c",x"40",x"40",x"7c"),
  2049 => (x"1c",x"00",x"00",x"7c"),
  2050 => (x"3c",x"60",x"60",x"3c"),
  2051 => (x"7c",x"3c",x"00",x"1c"),
  2052 => (x"7c",x"60",x"30",x"60"),
  2053 => (x"6c",x"44",x"00",x"3c"),
  2054 => (x"6c",x"38",x"10",x"38"),
  2055 => (x"1c",x"00",x"00",x"44"),
  2056 => (x"3c",x"60",x"e0",x"bc"),
  2057 => (x"44",x"00",x"00",x"1c"),
  2058 => (x"4c",x"5c",x"74",x"64"),
  2059 => (x"08",x"00",x"00",x"44"),
  2060 => (x"41",x"77",x"3e",x"08"),
  2061 => (x"00",x"00",x"00",x"41"),
  2062 => (x"00",x"7f",x"7f",x"00"),
  2063 => (x"41",x"00",x"00",x"00"),
  2064 => (x"08",x"3e",x"77",x"41"),
  2065 => (x"01",x"02",x"00",x"08"),
  2066 => (x"02",x"02",x"03",x"01"),
  2067 => (x"7f",x"7f",x"00",x"01"),
  2068 => (x"7f",x"7f",x"7f",x"7f"),
  2069 => (x"08",x"08",x"00",x"7f"),
  2070 => (x"3e",x"3e",x"1c",x"1c"),
  2071 => (x"7f",x"7f",x"7f",x"7f"),
  2072 => (x"1c",x"1c",x"3e",x"3e"),
  2073 => (x"10",x"00",x"08",x"08"),
  2074 => (x"18",x"7c",x"7c",x"18"),
  2075 => (x"10",x"00",x"00",x"10"),
  2076 => (x"30",x"7c",x"7c",x"30"),
  2077 => (x"30",x"10",x"00",x"10"),
  2078 => (x"1e",x"78",x"60",x"60"),
  2079 => (x"66",x"42",x"00",x"06"),
  2080 => (x"66",x"3c",x"18",x"3c"),
  2081 => (x"38",x"78",x"00",x"42"),
  2082 => (x"6c",x"c6",x"c2",x"6a"),
  2083 => (x"00",x"60",x"00",x"38"),
  2084 => (x"00",x"00",x"60",x"00"),
  2085 => (x"5e",x"0e",x"00",x"60"),
  2086 => (x"0e",x"5d",x"5c",x"5b"),
  2087 => (x"c2",x"4c",x"71",x"1e"),
  2088 => (x"4d",x"bf",x"d9",x"ee"),
  2089 => (x"1e",x"c0",x"4b",x"c0"),
  2090 => (x"c7",x"02",x"ab",x"74"),
  2091 => (x"48",x"a6",x"c4",x"87"),
  2092 => (x"87",x"c5",x"78",x"c0"),
  2093 => (x"c1",x"48",x"a6",x"c4"),
  2094 => (x"1e",x"66",x"c4",x"78"),
  2095 => (x"df",x"ee",x"49",x"73"),
  2096 => (x"c0",x"86",x"c8",x"87"),
  2097 => (x"ee",x"ef",x"49",x"e0"),
  2098 => (x"4a",x"a5",x"c4",x"87"),
  2099 => (x"f0",x"f0",x"49",x"6a"),
  2100 => (x"87",x"c6",x"f1",x"87"),
  2101 => (x"83",x"c1",x"85",x"cb"),
  2102 => (x"04",x"ab",x"b7",x"c8"),
  2103 => (x"26",x"87",x"c7",x"ff"),
  2104 => (x"4c",x"26",x"4d",x"26"),
  2105 => (x"4f",x"26",x"4b",x"26"),
  2106 => (x"c2",x"4a",x"71",x"1e"),
  2107 => (x"c2",x"5a",x"dd",x"ee"),
  2108 => (x"c7",x"48",x"dd",x"ee"),
  2109 => (x"dd",x"fe",x"49",x"78"),
  2110 => (x"1e",x"4f",x"26",x"87"),
  2111 => (x"4a",x"71",x"1e",x"73"),
  2112 => (x"03",x"aa",x"b7",x"c0"),
  2113 => (x"d2",x"c2",x"87",x"d3"),
  2114 => (x"c4",x"05",x"bf",x"fe"),
  2115 => (x"c2",x"4b",x"c1",x"87"),
  2116 => (x"c2",x"4b",x"c0",x"87"),
  2117 => (x"c4",x"5b",x"c2",x"d3"),
  2118 => (x"c2",x"d3",x"c2",x"87"),
  2119 => (x"fe",x"d2",x"c2",x"5a"),
  2120 => (x"9a",x"c1",x"4a",x"bf"),
  2121 => (x"49",x"a2",x"c0",x"c1"),
  2122 => (x"fc",x"87",x"e8",x"ec"),
  2123 => (x"fe",x"d2",x"c2",x"48"),
  2124 => (x"ef",x"fe",x"78",x"bf"),
  2125 => (x"4a",x"71",x"1e",x"87"),
  2126 => (x"72",x"1e",x"66",x"c4"),
  2127 => (x"87",x"f9",x"ea",x"49"),
  2128 => (x"1e",x"4f",x"26",x"26"),
  2129 => (x"c3",x"48",x"d4",x"ff"),
  2130 => (x"d0",x"ff",x"78",x"ff"),
  2131 => (x"78",x"e1",x"c0",x"48"),
  2132 => (x"c1",x"48",x"d4",x"ff"),
  2133 => (x"c4",x"48",x"71",x"78"),
  2134 => (x"08",x"d4",x"ff",x"30"),
  2135 => (x"48",x"d0",x"ff",x"78"),
  2136 => (x"26",x"78",x"e0",x"c0"),
  2137 => (x"d2",x"c2",x"1e",x"4f"),
  2138 => (x"e6",x"49",x"bf",x"fe"),
  2139 => (x"ee",x"c2",x"87",x"f9"),
  2140 => (x"bf",x"e8",x"48",x"d1"),
  2141 => (x"cd",x"ee",x"c2",x"78"),
  2142 => (x"78",x"bf",x"ec",x"48"),
  2143 => (x"bf",x"d1",x"ee",x"c2"),
  2144 => (x"ff",x"c3",x"49",x"4a"),
  2145 => (x"2a",x"b7",x"c8",x"99"),
  2146 => (x"b0",x"71",x"48",x"72"),
  2147 => (x"58",x"d9",x"ee",x"c2"),
  2148 => (x"5e",x"0e",x"4f",x"26"),
  2149 => (x"0e",x"5d",x"5c",x"5b"),
  2150 => (x"c8",x"ff",x"4b",x"71"),
  2151 => (x"cc",x"ee",x"c2",x"87"),
  2152 => (x"73",x"50",x"c0",x"48"),
  2153 => (x"87",x"df",x"e6",x"49"),
  2154 => (x"c2",x"4c",x"49",x"70"),
  2155 => (x"49",x"ee",x"cb",x"9c"),
  2156 => (x"70",x"87",x"d3",x"cc"),
  2157 => (x"cc",x"ee",x"c2",x"4d"),
  2158 => (x"c1",x"05",x"bf",x"97"),
  2159 => (x"66",x"d0",x"87",x"e2"),
  2160 => (x"d5",x"ee",x"c2",x"49"),
  2161 => (x"d6",x"05",x"99",x"bf"),
  2162 => (x"49",x"66",x"d4",x"87"),
  2163 => (x"bf",x"cd",x"ee",x"c2"),
  2164 => (x"87",x"cb",x"05",x"99"),
  2165 => (x"ee",x"e5",x"49",x"73"),
  2166 => (x"02",x"98",x"70",x"87"),
  2167 => (x"c1",x"87",x"c1",x"c1"),
  2168 => (x"87",x"c1",x"fe",x"4c"),
  2169 => (x"e9",x"cb",x"49",x"75"),
  2170 => (x"02",x"98",x"70",x"87"),
  2171 => (x"ee",x"c2",x"87",x"c6"),
  2172 => (x"50",x"c1",x"48",x"cc"),
  2173 => (x"97",x"cc",x"ee",x"c2"),
  2174 => (x"e3",x"c0",x"05",x"bf"),
  2175 => (x"d5",x"ee",x"c2",x"87"),
  2176 => (x"66",x"d0",x"49",x"bf"),
  2177 => (x"d6",x"ff",x"05",x"99"),
  2178 => (x"cd",x"ee",x"c2",x"87"),
  2179 => (x"66",x"d4",x"49",x"bf"),
  2180 => (x"ca",x"ff",x"05",x"99"),
  2181 => (x"e4",x"49",x"73",x"87"),
  2182 => (x"98",x"70",x"87",x"ed"),
  2183 => (x"87",x"ff",x"fe",x"05"),
  2184 => (x"fb",x"fa",x"48",x"74"),
  2185 => (x"5b",x"5e",x"0e",x"87"),
  2186 => (x"f8",x"0e",x"5d",x"5c"),
  2187 => (x"4c",x"4d",x"c0",x"86"),
  2188 => (x"c4",x"7e",x"bf",x"ec"),
  2189 => (x"ee",x"c2",x"48",x"a6"),
  2190 => (x"c1",x"78",x"bf",x"d9"),
  2191 => (x"c7",x"1e",x"c0",x"1e"),
  2192 => (x"87",x"ce",x"fd",x"49"),
  2193 => (x"98",x"70",x"86",x"c8"),
  2194 => (x"ff",x"87",x"cd",x"02"),
  2195 => (x"87",x"eb",x"fa",x"49"),
  2196 => (x"e3",x"49",x"da",x"c1"),
  2197 => (x"4d",x"c1",x"87",x"f1"),
  2198 => (x"97",x"cc",x"ee",x"c2"),
  2199 => (x"87",x"cf",x"02",x"bf"),
  2200 => (x"bf",x"e6",x"d2",x"c2"),
  2201 => (x"c2",x"b9",x"c1",x"49"),
  2202 => (x"71",x"59",x"ea",x"d2"),
  2203 => (x"c2",x"87",x"d4",x"fb"),
  2204 => (x"4b",x"bf",x"d1",x"ee"),
  2205 => (x"bf",x"fe",x"d2",x"c2"),
  2206 => (x"87",x"d9",x"c1",x"05"),
  2207 => (x"c8",x"48",x"a6",x"c4"),
  2208 => (x"c2",x"78",x"c0",x"c0"),
  2209 => (x"6e",x"7e",x"ea",x"d2"),
  2210 => (x"6e",x"49",x"bf",x"97"),
  2211 => (x"70",x"80",x"c1",x"48"),
  2212 => (x"f2",x"e2",x"71",x"7e"),
  2213 => (x"02",x"98",x"70",x"87"),
  2214 => (x"66",x"c4",x"87",x"c3"),
  2215 => (x"48",x"66",x"c4",x"b3"),
  2216 => (x"c8",x"28",x"b7",x"c1"),
  2217 => (x"98",x"70",x"58",x"a6"),
  2218 => (x"87",x"db",x"ff",x"05"),
  2219 => (x"e2",x"49",x"fd",x"c3"),
  2220 => (x"fa",x"c3",x"87",x"d5"),
  2221 => (x"87",x"cf",x"e2",x"49"),
  2222 => (x"ff",x"c3",x"49",x"73"),
  2223 => (x"c0",x"1e",x"71",x"99"),
  2224 => (x"87",x"f1",x"f9",x"49"),
  2225 => (x"b7",x"c8",x"49",x"73"),
  2226 => (x"c1",x"1e",x"71",x"29"),
  2227 => (x"87",x"e5",x"f9",x"49"),
  2228 => (x"fa",x"c5",x"86",x"c8"),
  2229 => (x"d5",x"ee",x"c2",x"87"),
  2230 => (x"02",x"9b",x"4b",x"bf"),
  2231 => (x"d2",x"c2",x"87",x"dd"),
  2232 => (x"c7",x"49",x"bf",x"fa"),
  2233 => (x"98",x"70",x"87",x"ec"),
  2234 => (x"c0",x"87",x"c4",x"05"),
  2235 => (x"c2",x"87",x"d2",x"4b"),
  2236 => (x"d1",x"c7",x"49",x"e0"),
  2237 => (x"fe",x"d2",x"c2",x"87"),
  2238 => (x"c2",x"87",x"c6",x"58"),
  2239 => (x"c0",x"48",x"fa",x"d2"),
  2240 => (x"c2",x"49",x"73",x"78"),
  2241 => (x"87",x"ce",x"05",x"99"),
  2242 => (x"e0",x"49",x"eb",x"c3"),
  2243 => (x"49",x"70",x"87",x"f9"),
  2244 => (x"c0",x"02",x"99",x"c2"),
  2245 => (x"4c",x"fb",x"87",x"c2"),
  2246 => (x"99",x"c1",x"49",x"73"),
  2247 => (x"c3",x"87",x"ce",x"05"),
  2248 => (x"e2",x"e0",x"49",x"f4"),
  2249 => (x"c2",x"49",x"70",x"87"),
  2250 => (x"c2",x"c0",x"02",x"99"),
  2251 => (x"73",x"4c",x"fa",x"87"),
  2252 => (x"05",x"99",x"c8",x"49"),
  2253 => (x"f5",x"c3",x"87",x"cd"),
  2254 => (x"87",x"cb",x"e0",x"49"),
  2255 => (x"99",x"c2",x"49",x"70"),
  2256 => (x"c2",x"87",x"d6",x"02"),
  2257 => (x"02",x"bf",x"dd",x"ee"),
  2258 => (x"48",x"87",x"ca",x"c0"),
  2259 => (x"ee",x"c2",x"88",x"c1"),
  2260 => (x"c2",x"c0",x"58",x"e1"),
  2261 => (x"c1",x"4c",x"ff",x"87"),
  2262 => (x"c4",x"49",x"73",x"4d"),
  2263 => (x"ce",x"c0",x"05",x"99"),
  2264 => (x"49",x"f2",x"c3",x"87"),
  2265 => (x"87",x"df",x"df",x"ff"),
  2266 => (x"99",x"c2",x"49",x"70"),
  2267 => (x"c2",x"87",x"dc",x"02"),
  2268 => (x"7e",x"bf",x"dd",x"ee"),
  2269 => (x"a8",x"b7",x"c7",x"48"),
  2270 => (x"87",x"cb",x"c0",x"03"),
  2271 => (x"80",x"c1",x"48",x"6e"),
  2272 => (x"58",x"e1",x"ee",x"c2"),
  2273 => (x"fe",x"87",x"c2",x"c0"),
  2274 => (x"c3",x"4d",x"c1",x"4c"),
  2275 => (x"de",x"ff",x"49",x"fd"),
  2276 => (x"49",x"70",x"87",x"f5"),
  2277 => (x"c0",x"02",x"99",x"c2"),
  2278 => (x"ee",x"c2",x"87",x"d5"),
  2279 => (x"c0",x"02",x"bf",x"dd"),
  2280 => (x"ee",x"c2",x"87",x"c9"),
  2281 => (x"78",x"c0",x"48",x"dd"),
  2282 => (x"fd",x"87",x"c2",x"c0"),
  2283 => (x"c3",x"4d",x"c1",x"4c"),
  2284 => (x"de",x"ff",x"49",x"fa"),
  2285 => (x"49",x"70",x"87",x"d1"),
  2286 => (x"c0",x"02",x"99",x"c2"),
  2287 => (x"ee",x"c2",x"87",x"d9"),
  2288 => (x"c7",x"48",x"bf",x"dd"),
  2289 => (x"c0",x"03",x"a8",x"b7"),
  2290 => (x"ee",x"c2",x"87",x"c9"),
  2291 => (x"78",x"c7",x"48",x"dd"),
  2292 => (x"fc",x"87",x"c2",x"c0"),
  2293 => (x"c0",x"4d",x"c1",x"4c"),
  2294 => (x"c0",x"03",x"ac",x"b7"),
  2295 => (x"66",x"c4",x"87",x"d3"),
  2296 => (x"80",x"d8",x"c1",x"48"),
  2297 => (x"bf",x"6e",x"7e",x"70"),
  2298 => (x"87",x"c5",x"c0",x"02"),
  2299 => (x"73",x"49",x"74",x"4b"),
  2300 => (x"c3",x"1e",x"c0",x"0f"),
  2301 => (x"da",x"c1",x"1e",x"f0"),
  2302 => (x"87",x"d6",x"f6",x"49"),
  2303 => (x"98",x"70",x"86",x"c8"),
  2304 => (x"87",x"d8",x"c0",x"02"),
  2305 => (x"bf",x"dd",x"ee",x"c2"),
  2306 => (x"cb",x"49",x"6e",x"7e"),
  2307 => (x"4a",x"66",x"c4",x"91"),
  2308 => (x"02",x"6a",x"82",x"71"),
  2309 => (x"4b",x"87",x"c5",x"c0"),
  2310 => (x"0f",x"73",x"49",x"6e"),
  2311 => (x"c0",x"02",x"9d",x"75"),
  2312 => (x"ee",x"c2",x"87",x"c8"),
  2313 => (x"f1",x"49",x"bf",x"dd"),
  2314 => (x"d3",x"c2",x"87",x"ec"),
  2315 => (x"c0",x"02",x"bf",x"c2"),
  2316 => (x"c2",x"49",x"87",x"dd"),
  2317 => (x"98",x"70",x"87",x"dc"),
  2318 => (x"87",x"d3",x"c0",x"02"),
  2319 => (x"bf",x"dd",x"ee",x"c2"),
  2320 => (x"87",x"d2",x"f1",x"49"),
  2321 => (x"f2",x"f2",x"49",x"c0"),
  2322 => (x"c2",x"d3",x"c2",x"87"),
  2323 => (x"f8",x"78",x"c0",x"48"),
  2324 => (x"87",x"cc",x"f2",x"8e"),
  2325 => (x"5c",x"5b",x"5e",x"0e"),
  2326 => (x"71",x"1e",x"0e",x"5d"),
  2327 => (x"d9",x"ee",x"c2",x"4c"),
  2328 => (x"cd",x"c1",x"49",x"bf"),
  2329 => (x"d1",x"c1",x"4d",x"a1"),
  2330 => (x"74",x"7e",x"69",x"81"),
  2331 => (x"87",x"cf",x"02",x"9c"),
  2332 => (x"74",x"4b",x"a5",x"c4"),
  2333 => (x"d9",x"ee",x"c2",x"7b"),
  2334 => (x"eb",x"f1",x"49",x"bf"),
  2335 => (x"74",x"7b",x"6e",x"87"),
  2336 => (x"87",x"c4",x"05",x"9c"),
  2337 => (x"87",x"c2",x"4b",x"c0"),
  2338 => (x"49",x"73",x"4b",x"c1"),
  2339 => (x"d4",x"87",x"ec",x"f1"),
  2340 => (x"87",x"c8",x"02",x"66"),
  2341 => (x"87",x"ee",x"c0",x"49"),
  2342 => (x"87",x"c2",x"4a",x"70"),
  2343 => (x"d3",x"c2",x"4a",x"c0"),
  2344 => (x"f0",x"26",x"5a",x"c6"),
  2345 => (x"00",x"00",x"87",x"fa"),
  2346 => (x"12",x"58",x"00",x"00"),
  2347 => (x"1b",x"1d",x"14",x"11"),
  2348 => (x"59",x"5a",x"23",x"1c"),
  2349 => (x"f2",x"f5",x"94",x"91"),
  2350 => (x"00",x"00",x"f4",x"eb"),
  2351 => (x"00",x"00",x"00",x"00"),
  2352 => (x"00",x"00",x"00",x"00"),
  2353 => (x"71",x"1e",x"00",x"00"),
  2354 => (x"bf",x"c8",x"ff",x"4a"),
  2355 => (x"48",x"a1",x"72",x"49"),
  2356 => (x"ff",x"1e",x"4f",x"26"),
  2357 => (x"fe",x"89",x"bf",x"c8"),
  2358 => (x"c0",x"c0",x"c0",x"c0"),
  2359 => (x"c4",x"01",x"a9",x"c0"),
  2360 => (x"c2",x"4a",x"c0",x"87"),
  2361 => (x"72",x"4a",x"c1",x"87"),
  2362 => (x"0e",x"4f",x"26",x"48"),
  2363 => (x"5d",x"5c",x"5b",x"5e"),
  2364 => (x"ff",x"4b",x"71",x"0e"),
  2365 => (x"66",x"d0",x"4c",x"d4"),
  2366 => (x"d6",x"78",x"c0",x"48"),
  2367 => (x"fe",x"da",x"ff",x"49"),
  2368 => (x"7c",x"ff",x"c3",x"87"),
  2369 => (x"ff",x"c3",x"49",x"6c"),
  2370 => (x"49",x"4d",x"71",x"99"),
  2371 => (x"c1",x"99",x"f0",x"c3"),
  2372 => (x"cb",x"05",x"a9",x"e0"),
  2373 => (x"7c",x"ff",x"c3",x"87"),
  2374 => (x"98",x"c3",x"48",x"6c"),
  2375 => (x"78",x"08",x"66",x"d0"),
  2376 => (x"6c",x"7c",x"ff",x"c3"),
  2377 => (x"31",x"c8",x"49",x"4a"),
  2378 => (x"6c",x"7c",x"ff",x"c3"),
  2379 => (x"72",x"b2",x"71",x"4a"),
  2380 => (x"c3",x"31",x"c8",x"49"),
  2381 => (x"4a",x"6c",x"7c",x"ff"),
  2382 => (x"49",x"72",x"b2",x"71"),
  2383 => (x"ff",x"c3",x"31",x"c8"),
  2384 => (x"71",x"4a",x"6c",x"7c"),
  2385 => (x"48",x"d0",x"ff",x"b2"),
  2386 => (x"73",x"78",x"e0",x"c0"),
  2387 => (x"87",x"c2",x"02",x"9b"),
  2388 => (x"48",x"75",x"7b",x"72"),
  2389 => (x"4c",x"26",x"4d",x"26"),
  2390 => (x"4f",x"26",x"4b",x"26"),
  2391 => (x"0e",x"4f",x"26",x"1e"),
  2392 => (x"0e",x"5c",x"5b",x"5e"),
  2393 => (x"1e",x"76",x"86",x"f8"),
  2394 => (x"fd",x"49",x"a6",x"c8"),
  2395 => (x"86",x"c4",x"87",x"fd"),
  2396 => (x"48",x"6e",x"4b",x"70"),
  2397 => (x"c2",x"03",x"a8",x"c2"),
  2398 => (x"4a",x"73",x"87",x"f0"),
  2399 => (x"c1",x"9a",x"f0",x"c3"),
  2400 => (x"c7",x"02",x"aa",x"d0"),
  2401 => (x"aa",x"e0",x"c1",x"87"),
  2402 => (x"87",x"de",x"c2",x"05"),
  2403 => (x"99",x"c8",x"49",x"73"),
  2404 => (x"ff",x"87",x"c3",x"02"),
  2405 => (x"4c",x"73",x"87",x"c6"),
  2406 => (x"ac",x"c2",x"9c",x"c3"),
  2407 => (x"87",x"c2",x"c1",x"05"),
  2408 => (x"c9",x"49",x"66",x"c4"),
  2409 => (x"c4",x"1e",x"71",x"31"),
  2410 => (x"92",x"d4",x"4a",x"66"),
  2411 => (x"49",x"e1",x"ee",x"c2"),
  2412 => (x"d0",x"fe",x"81",x"72"),
  2413 => (x"49",x"d8",x"87",x"d1"),
  2414 => (x"87",x"c3",x"d8",x"ff"),
  2415 => (x"c2",x"1e",x"c0",x"c8"),
  2416 => (x"fd",x"49",x"fe",x"dc"),
  2417 => (x"ff",x"87",x"d7",x"ec"),
  2418 => (x"e0",x"c0",x"48",x"d0"),
  2419 => (x"fe",x"dc",x"c2",x"78"),
  2420 => (x"4a",x"66",x"cc",x"1e"),
  2421 => (x"ee",x"c2",x"92",x"d4"),
  2422 => (x"81",x"72",x"49",x"e1"),
  2423 => (x"87",x"d9",x"ce",x"fe"),
  2424 => (x"ac",x"c1",x"86",x"cc"),
  2425 => (x"87",x"c2",x"c1",x"05"),
  2426 => (x"c9",x"49",x"66",x"c4"),
  2427 => (x"c4",x"1e",x"71",x"31"),
  2428 => (x"92",x"d4",x"4a",x"66"),
  2429 => (x"49",x"e1",x"ee",x"c2"),
  2430 => (x"cf",x"fe",x"81",x"72"),
  2431 => (x"dc",x"c2",x"87",x"c9"),
  2432 => (x"66",x"c8",x"1e",x"fe"),
  2433 => (x"c2",x"92",x"d4",x"4a"),
  2434 => (x"72",x"49",x"e1",x"ee"),
  2435 => (x"da",x"cc",x"fe",x"81"),
  2436 => (x"ff",x"49",x"d7",x"87"),
  2437 => (x"c8",x"87",x"e8",x"d6"),
  2438 => (x"dc",x"c2",x"1e",x"c0"),
  2439 => (x"ea",x"fd",x"49",x"fe"),
  2440 => (x"86",x"cc",x"87",x"d5"),
  2441 => (x"c0",x"48",x"d0",x"ff"),
  2442 => (x"8e",x"f8",x"78",x"e0"),
  2443 => (x"0e",x"87",x"e7",x"fc"),
  2444 => (x"5d",x"5c",x"5b",x"5e"),
  2445 => (x"4d",x"71",x"1e",x"0e"),
  2446 => (x"d4",x"4c",x"d4",x"ff"),
  2447 => (x"c3",x"48",x"7e",x"66"),
  2448 => (x"c5",x"06",x"a8",x"b7"),
  2449 => (x"c1",x"48",x"c0",x"87"),
  2450 => (x"49",x"75",x"87",x"e9"),
  2451 => (x"87",x"ff",x"dc",x"fe"),
  2452 => (x"66",x"c4",x"1e",x"75"),
  2453 => (x"c2",x"93",x"d4",x"4b"),
  2454 => (x"73",x"83",x"e1",x"ee"),
  2455 => (x"d8",x"c6",x"fe",x"49"),
  2456 => (x"6b",x"83",x"c8",x"87"),
  2457 => (x"48",x"d0",x"ff",x"4b"),
  2458 => (x"dd",x"78",x"e1",x"c8"),
  2459 => (x"c3",x"48",x"73",x"7c"),
  2460 => (x"7c",x"70",x"98",x"ff"),
  2461 => (x"b7",x"c8",x"49",x"73"),
  2462 => (x"c3",x"48",x"71",x"29"),
  2463 => (x"7c",x"70",x"98",x"ff"),
  2464 => (x"b7",x"d0",x"49",x"73"),
  2465 => (x"c3",x"48",x"71",x"29"),
  2466 => (x"7c",x"70",x"98",x"ff"),
  2467 => (x"b7",x"d8",x"48",x"73"),
  2468 => (x"c0",x"7c",x"70",x"28"),
  2469 => (x"7c",x"7c",x"7c",x"7c"),
  2470 => (x"7c",x"7c",x"7c",x"7c"),
  2471 => (x"7c",x"7c",x"7c",x"7c"),
  2472 => (x"c0",x"48",x"d0",x"ff"),
  2473 => (x"66",x"c4",x"78",x"e0"),
  2474 => (x"ff",x"49",x"dc",x"1e"),
  2475 => (x"c8",x"87",x"f5",x"d4"),
  2476 => (x"26",x"48",x"73",x"86"),
  2477 => (x"1e",x"87",x"dd",x"fa"),
  2478 => (x"4b",x"c0",x"1e",x"73"),
  2479 => (x"f8",x"db",x"c2",x"1e"),
  2480 => (x"ea",x"fd",x"49",x"bf"),
  2481 => (x"c2",x"86",x"c4",x"87"),
  2482 => (x"49",x"bf",x"fc",x"db"),
  2483 => (x"87",x"e3",x"de",x"fe"),
  2484 => (x"c4",x"05",x"98",x"70"),
  2485 => (x"e5",x"db",x"c2",x"87"),
  2486 => (x"c4",x"48",x"73",x"4b"),
  2487 => (x"26",x"4d",x"26",x"87"),
  2488 => (x"26",x"4b",x"26",x"4c"),
  2489 => (x"4d",x"4f",x"52",x"4f"),
  2490 => (x"61",x"6f",x"6c",x"20"),
  2491 => (x"67",x"6e",x"69",x"64"),
  2492 => (x"69",x"61",x"66",x"20"),
  2493 => (x"00",x"64",x"65",x"6c"),
  2494 => (x"00",x"00",x"27",x"00"),
  2495 => (x"00",x"00",x"27",x"0c"),
  2496 => (x"20",x"43",x"42",x"42"),
  2497 => (x"20",x"20",x"20",x"20"),
  2498 => (x"00",x"44",x"48",x"56"),
  2499 => (x"20",x"43",x"42",x"42"),
  2500 => (x"20",x"20",x"20",x"20"),
  2501 => (x"00",x"4d",x"4f",x"52"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

