
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"3e",x"7f",x"4d"),
     1 => (x"7f",x"06",x"04",x"00"),
     2 => (x"00",x"00",x"00",x"7f"),
     3 => (x"71",x"63",x"42",x"00"),
     4 => (x"00",x"46",x"4f",x"59"),
     5 => (x"49",x"63",x"22",x"00"),
     6 => (x"00",x"36",x"7f",x"49"),
     7 => (x"13",x"16",x"1c",x"18"),
     8 => (x"00",x"10",x"7f",x"7f"),
     9 => (x"45",x"67",x"27",x"00"),
    10 => (x"00",x"39",x"7d",x"45"),
    11 => (x"4b",x"7e",x"3c",x"00"),
    12 => (x"00",x"30",x"79",x"49"),
    13 => (x"71",x"01",x"01",x"00"),
    14 => (x"00",x"07",x"0f",x"79"),
    15 => (x"49",x"7f",x"36",x"00"),
    16 => (x"00",x"36",x"7f",x"49"),
    17 => (x"49",x"4f",x"06",x"00"),
    18 => (x"00",x"1e",x"3f",x"69"),
    19 => (x"66",x"00",x"00",x"00"),
    20 => (x"00",x"00",x"00",x"66"),
    21 => (x"e6",x"80",x"00",x"00"),
    22 => (x"00",x"00",x"00",x"66"),
    23 => (x"14",x"08",x"08",x"00"),
    24 => (x"00",x"22",x"22",x"14"),
    25 => (x"14",x"14",x"14",x"00"),
    26 => (x"00",x"14",x"14",x"14"),
    27 => (x"14",x"22",x"22",x"00"),
    28 => (x"00",x"08",x"08",x"14"),
    29 => (x"51",x"03",x"02",x"00"),
    30 => (x"00",x"06",x"0f",x"59"),
    31 => (x"5d",x"41",x"7f",x"3e"),
    32 => (x"00",x"1e",x"1f",x"55"),
    33 => (x"09",x"7f",x"7e",x"00"),
    34 => (x"00",x"7e",x"7f",x"09"),
    35 => (x"49",x"7f",x"7f",x"00"),
    36 => (x"00",x"36",x"7f",x"49"),
    37 => (x"63",x"3e",x"1c",x"00"),
    38 => (x"00",x"41",x"41",x"41"),
    39 => (x"41",x"7f",x"7f",x"00"),
    40 => (x"00",x"1c",x"3e",x"63"),
    41 => (x"49",x"7f",x"7f",x"00"),
    42 => (x"00",x"41",x"41",x"49"),
    43 => (x"09",x"7f",x"7f",x"00"),
    44 => (x"00",x"01",x"01",x"09"),
    45 => (x"41",x"7f",x"3e",x"00"),
    46 => (x"00",x"7a",x"7b",x"49"),
    47 => (x"08",x"7f",x"7f",x"00"),
    48 => (x"00",x"7f",x"7f",x"08"),
    49 => (x"7f",x"41",x"00",x"00"),
    50 => (x"00",x"00",x"41",x"7f"),
    51 => (x"40",x"60",x"20",x"00"),
    52 => (x"00",x"3f",x"7f",x"40"),
    53 => (x"1c",x"08",x"7f",x"7f"),
    54 => (x"00",x"41",x"63",x"36"),
    55 => (x"40",x"7f",x"7f",x"00"),
    56 => (x"00",x"40",x"40",x"40"),
    57 => (x"0c",x"06",x"7f",x"7f"),
    58 => (x"00",x"7f",x"7f",x"06"),
    59 => (x"0c",x"06",x"7f",x"7f"),
    60 => (x"00",x"7f",x"7f",x"18"),
    61 => (x"41",x"7f",x"3e",x"00"),
    62 => (x"00",x"3e",x"7f",x"41"),
    63 => (x"09",x"7f",x"7f",x"00"),
    64 => (x"00",x"06",x"0f",x"09"),
    65 => (x"61",x"41",x"7f",x"3e"),
    66 => (x"00",x"40",x"7e",x"7f"),
    67 => (x"09",x"7f",x"7f",x"00"),
    68 => (x"00",x"66",x"7f",x"19"),
    69 => (x"4d",x"6f",x"26",x"00"),
    70 => (x"00",x"32",x"7b",x"59"),
    71 => (x"7f",x"01",x"01",x"00"),
    72 => (x"00",x"01",x"01",x"7f"),
    73 => (x"40",x"7f",x"3f",x"00"),
    74 => (x"00",x"3f",x"7f",x"40"),
    75 => (x"70",x"3f",x"0f",x"00"),
    76 => (x"00",x"0f",x"3f",x"70"),
    77 => (x"18",x"30",x"7f",x"7f"),
    78 => (x"00",x"7f",x"7f",x"30"),
    79 => (x"1c",x"36",x"63",x"41"),
    80 => (x"41",x"63",x"36",x"1c"),
    81 => (x"7c",x"06",x"03",x"01"),
    82 => (x"01",x"03",x"06",x"7c"),
    83 => (x"4d",x"59",x"71",x"61"),
    84 => (x"00",x"41",x"43",x"47"),
    85 => (x"7f",x"7f",x"00",x"00"),
    86 => (x"00",x"00",x"41",x"41"),
    87 => (x"0c",x"06",x"03",x"01"),
    88 => (x"40",x"60",x"30",x"18"),
    89 => (x"41",x"41",x"00",x"00"),
    90 => (x"00",x"00",x"7f",x"7f"),
    91 => (x"03",x"06",x"0c",x"08"),
    92 => (x"00",x"08",x"0c",x"06"),
    93 => (x"80",x"80",x"80",x"80"),
    94 => (x"00",x"80",x"80",x"80"),
    95 => (x"03",x"00",x"00",x"00"),
    96 => (x"00",x"00",x"04",x"07"),
    97 => (x"54",x"74",x"20",x"00"),
    98 => (x"00",x"78",x"7c",x"54"),
    99 => (x"44",x"7f",x"7f",x"00"),
   100 => (x"00",x"38",x"7c",x"44"),
   101 => (x"44",x"7c",x"38",x"00"),
   102 => (x"00",x"00",x"44",x"44"),
   103 => (x"44",x"7c",x"38",x"00"),
   104 => (x"00",x"7f",x"7f",x"44"),
   105 => (x"54",x"7c",x"38",x"00"),
   106 => (x"00",x"18",x"5c",x"54"),
   107 => (x"7f",x"7e",x"04",x"00"),
   108 => (x"00",x"00",x"05",x"05"),
   109 => (x"a4",x"bc",x"18",x"00"),
   110 => (x"00",x"7c",x"fc",x"a4"),
   111 => (x"04",x"7f",x"7f",x"00"),
   112 => (x"00",x"78",x"7c",x"04"),
   113 => (x"3d",x"00",x"00",x"00"),
   114 => (x"00",x"00",x"40",x"7d"),
   115 => (x"80",x"80",x"80",x"00"),
   116 => (x"00",x"00",x"7d",x"fd"),
   117 => (x"10",x"7f",x"7f",x"00"),
   118 => (x"00",x"44",x"6c",x"38"),
   119 => (x"3f",x"00",x"00",x"00"),
   120 => (x"00",x"00",x"40",x"7f"),
   121 => (x"18",x"0c",x"7c",x"7c"),
   122 => (x"00",x"78",x"7c",x"0c"),
   123 => (x"04",x"7c",x"7c",x"00"),
   124 => (x"00",x"78",x"7c",x"04"),
   125 => (x"44",x"7c",x"38",x"00"),
   126 => (x"00",x"38",x"7c",x"44"),
   127 => (x"24",x"fc",x"fc",x"00"),
   128 => (x"00",x"18",x"3c",x"24"),
   129 => (x"24",x"3c",x"18",x"00"),
   130 => (x"00",x"fc",x"fc",x"24"),
   131 => (x"04",x"7c",x"7c",x"00"),
   132 => (x"00",x"08",x"0c",x"04"),
   133 => (x"54",x"5c",x"48",x"00"),
   134 => (x"00",x"20",x"74",x"54"),
   135 => (x"7f",x"3f",x"04",x"00"),
   136 => (x"00",x"00",x"44",x"44"),
   137 => (x"40",x"7c",x"3c",x"00"),
   138 => (x"00",x"7c",x"7c",x"40"),
   139 => (x"60",x"3c",x"1c",x"00"),
   140 => (x"00",x"1c",x"3c",x"60"),
   141 => (x"30",x"60",x"7c",x"3c"),
   142 => (x"00",x"3c",x"7c",x"60"),
   143 => (x"10",x"38",x"6c",x"44"),
   144 => (x"00",x"44",x"6c",x"38"),
   145 => (x"e0",x"bc",x"1c",x"00"),
   146 => (x"00",x"1c",x"3c",x"60"),
   147 => (x"74",x"64",x"44",x"00"),
   148 => (x"00",x"44",x"4c",x"5c"),
   149 => (x"3e",x"08",x"08",x"00"),
   150 => (x"00",x"41",x"41",x"77"),
   151 => (x"7f",x"00",x"00",x"00"),
   152 => (x"00",x"00",x"00",x"7f"),
   153 => (x"77",x"41",x"41",x"00"),
   154 => (x"00",x"08",x"08",x"3e"),
   155 => (x"03",x"01",x"01",x"02"),
   156 => (x"00",x"01",x"02",x"02"),
   157 => (x"7f",x"7f",x"7f",x"7f"),
   158 => (x"00",x"7f",x"7f",x"7f"),
   159 => (x"1c",x"1c",x"08",x"08"),
   160 => (x"7f",x"7f",x"3e",x"3e"),
   161 => (x"3e",x"3e",x"7f",x"7f"),
   162 => (x"08",x"08",x"1c",x"1c"),
   163 => (x"7c",x"18",x"10",x"00"),
   164 => (x"00",x"10",x"18",x"7c"),
   165 => (x"7c",x"30",x"10",x"00"),
   166 => (x"00",x"10",x"30",x"7c"),
   167 => (x"60",x"60",x"30",x"10"),
   168 => (x"00",x"06",x"1e",x"78"),
   169 => (x"18",x"3c",x"66",x"42"),
   170 => (x"00",x"42",x"66",x"3c"),
   171 => (x"c2",x"6a",x"38",x"78"),
   172 => (x"00",x"38",x"6c",x"c6"),
   173 => (x"60",x"00",x"00",x"60"),
   174 => (x"00",x"60",x"00",x"00"),
   175 => (x"5c",x"5b",x"5e",x"0e"),
   176 => (x"86",x"fc",x"0e",x"5d"),
   177 => (x"f5",x"c2",x"7e",x"71"),
   178 => (x"c0",x"4c",x"bf",x"d4"),
   179 => (x"c4",x"1e",x"c0",x"4b"),
   180 => (x"c4",x"02",x"ab",x"66"),
   181 => (x"c2",x"4d",x"c0",x"87"),
   182 => (x"75",x"4d",x"c1",x"87"),
   183 => (x"ee",x"49",x"73",x"1e"),
   184 => (x"86",x"c8",x"87",x"e1"),
   185 => (x"ef",x"49",x"e0",x"c0"),
   186 => (x"a4",x"c4",x"87",x"ea"),
   187 => (x"f0",x"49",x"6a",x"4a"),
   188 => (x"c8",x"f1",x"87",x"f1"),
   189 => (x"c1",x"84",x"cc",x"87"),
   190 => (x"ab",x"b7",x"c8",x"83"),
   191 => (x"87",x"cd",x"ff",x"04"),
   192 => (x"4d",x"26",x"8e",x"fc"),
   193 => (x"4b",x"26",x"4c",x"26"),
   194 => (x"71",x"1e",x"4f",x"26"),
   195 => (x"d8",x"f5",x"c2",x"4a"),
   196 => (x"d8",x"f5",x"c2",x"5a"),
   197 => (x"49",x"78",x"c7",x"48"),
   198 => (x"26",x"87",x"e1",x"fe"),
   199 => (x"1e",x"73",x"1e",x"4f"),
   200 => (x"b7",x"c0",x"4a",x"71"),
   201 => (x"87",x"d3",x"03",x"aa"),
   202 => (x"bf",x"f8",x"d9",x"c2"),
   203 => (x"c1",x"87",x"c4",x"05"),
   204 => (x"c0",x"87",x"c2",x"4b"),
   205 => (x"fc",x"d9",x"c2",x"4b"),
   206 => (x"c2",x"87",x"c4",x"5b"),
   207 => (x"fc",x"5a",x"fc",x"d9"),
   208 => (x"f8",x"d9",x"c2",x"48"),
   209 => (x"c1",x"4a",x"78",x"bf"),
   210 => (x"a2",x"c0",x"c1",x"9a"),
   211 => (x"87",x"e6",x"ec",x"49"),
   212 => (x"4f",x"26",x"4b",x"26"),
   213 => (x"c4",x"4a",x"71",x"1e"),
   214 => (x"49",x"72",x"1e",x"66"),
   215 => (x"fc",x"87",x"f0",x"eb"),
   216 => (x"1e",x"4f",x"26",x"8e"),
   217 => (x"c3",x"48",x"d4",x"ff"),
   218 => (x"d0",x"ff",x"78",x"ff"),
   219 => (x"78",x"e1",x"c0",x"48"),
   220 => (x"c1",x"48",x"d4",x"ff"),
   221 => (x"c4",x"48",x"71",x"78"),
   222 => (x"08",x"d4",x"ff",x"30"),
   223 => (x"48",x"d0",x"ff",x"78"),
   224 => (x"26",x"78",x"e0",x"c0"),
   225 => (x"5b",x"5e",x"0e",x"4f"),
   226 => (x"ec",x"0e",x"5d",x"5c"),
   227 => (x"48",x"a6",x"c8",x"86"),
   228 => (x"c4",x"7e",x"78",x"c0"),
   229 => (x"78",x"bf",x"ec",x"80"),
   230 => (x"f5",x"c2",x"80",x"f8"),
   231 => (x"e8",x"78",x"bf",x"d4"),
   232 => (x"d9",x"c2",x"4c",x"bf"),
   233 => (x"e3",x"49",x"bf",x"f8"),
   234 => (x"ee",x"cb",x"87",x"eb"),
   235 => (x"87",x"cc",x"cb",x"49"),
   236 => (x"c7",x"58",x"a6",x"d4"),
   237 => (x"87",x"df",x"e7",x"49"),
   238 => (x"c9",x"05",x"98",x"70"),
   239 => (x"49",x"66",x"cc",x"87"),
   240 => (x"c1",x"02",x"99",x"c1"),
   241 => (x"66",x"d0",x"87",x"c4"),
   242 => (x"ec",x"7e",x"c1",x"4d"),
   243 => (x"d9",x"c2",x"4b",x"bf"),
   244 => (x"e2",x"49",x"bf",x"f8"),
   245 => (x"49",x"75",x"87",x"ff"),
   246 => (x"70",x"87",x"ed",x"ca"),
   247 => (x"87",x"d7",x"02",x"98"),
   248 => (x"bf",x"e0",x"d9",x"c2"),
   249 => (x"c2",x"b9",x"c1",x"49"),
   250 => (x"71",x"59",x"e4",x"d9"),
   251 => (x"cb",x"87",x"f4",x"fd"),
   252 => (x"c7",x"ca",x"49",x"ee"),
   253 => (x"c7",x"4d",x"70",x"87"),
   254 => (x"87",x"db",x"e6",x"49"),
   255 => (x"ff",x"05",x"98",x"70"),
   256 => (x"49",x"73",x"87",x"c7"),
   257 => (x"fe",x"05",x"99",x"c1"),
   258 => (x"02",x"6e",x"87",x"ff"),
   259 => (x"c2",x"87",x"e3",x"c0"),
   260 => (x"4a",x"bf",x"f8",x"d9"),
   261 => (x"d9",x"c2",x"ba",x"c1"),
   262 => (x"0a",x"fc",x"5a",x"fc"),
   263 => (x"9a",x"c1",x"0a",x"7a"),
   264 => (x"49",x"a2",x"c0",x"c1"),
   265 => (x"c1",x"87",x"cf",x"e9"),
   266 => (x"ea",x"e5",x"49",x"da"),
   267 => (x"48",x"a6",x"c8",x"87"),
   268 => (x"d9",x"c2",x"78",x"c1"),
   269 => (x"c1",x"05",x"bf",x"f8"),
   270 => (x"c0",x"c8",x"87",x"c5"),
   271 => (x"d9",x"c2",x"4d",x"c0"),
   272 => (x"49",x"13",x"4b",x"e4"),
   273 => (x"87",x"cf",x"e5",x"49"),
   274 => (x"c2",x"02",x"98",x"70"),
   275 => (x"c1",x"b4",x"75",x"87"),
   276 => (x"ff",x"05",x"2d",x"b7"),
   277 => (x"49",x"74",x"87",x"ec"),
   278 => (x"71",x"99",x"ff",x"c3"),
   279 => (x"fb",x"49",x"c0",x"1e"),
   280 => (x"49",x"74",x"87",x"f2"),
   281 => (x"71",x"29",x"b7",x"c8"),
   282 => (x"fb",x"49",x"c1",x"1e"),
   283 => (x"86",x"c8",x"87",x"e6"),
   284 => (x"e4",x"49",x"fd",x"c3"),
   285 => (x"fa",x"c3",x"87",x"e1"),
   286 => (x"87",x"db",x"e4",x"49"),
   287 => (x"74",x"87",x"d4",x"c7"),
   288 => (x"99",x"ff",x"c3",x"49"),
   289 => (x"71",x"2c",x"b7",x"c8"),
   290 => (x"02",x"9c",x"74",x"b4"),
   291 => (x"d9",x"c2",x"87",x"df"),
   292 => (x"c7",x"49",x"bf",x"f4"),
   293 => (x"98",x"70",x"87",x"f2"),
   294 => (x"87",x"c4",x"c0",x"05"),
   295 => (x"87",x"d3",x"4c",x"c0"),
   296 => (x"c7",x"49",x"e0",x"c2"),
   297 => (x"d9",x"c2",x"87",x"d6"),
   298 => (x"c6",x"c0",x"58",x"f8"),
   299 => (x"f4",x"d9",x"c2",x"87"),
   300 => (x"74",x"78",x"c0",x"48"),
   301 => (x"05",x"99",x"c8",x"49"),
   302 => (x"c3",x"87",x"ce",x"c0"),
   303 => (x"d6",x"e3",x"49",x"f5"),
   304 => (x"c2",x"49",x"70",x"87"),
   305 => (x"e7",x"c0",x"02",x"99"),
   306 => (x"d8",x"f5",x"c2",x"87"),
   307 => (x"ca",x"c0",x"02",x"bf"),
   308 => (x"88",x"c1",x"48",x"87"),
   309 => (x"58",x"dc",x"f5",x"c2"),
   310 => (x"c4",x"87",x"d0",x"c0"),
   311 => (x"e0",x"c1",x"4a",x"66"),
   312 => (x"c0",x"02",x"6a",x"82"),
   313 => (x"ff",x"4b",x"87",x"c5"),
   314 => (x"c8",x"0f",x"73",x"49"),
   315 => (x"78",x"c1",x"48",x"a6"),
   316 => (x"99",x"c4",x"49",x"74"),
   317 => (x"87",x"ce",x"c0",x"05"),
   318 => (x"e2",x"49",x"f2",x"c3"),
   319 => (x"49",x"70",x"87",x"d9"),
   320 => (x"c0",x"02",x"99",x"c2"),
   321 => (x"f5",x"c2",x"87",x"f0"),
   322 => (x"48",x"7e",x"bf",x"d8"),
   323 => (x"03",x"a8",x"b7",x"c7"),
   324 => (x"6e",x"87",x"cb",x"c0"),
   325 => (x"c2",x"80",x"c1",x"48"),
   326 => (x"c0",x"58",x"dc",x"f5"),
   327 => (x"66",x"c4",x"87",x"d3"),
   328 => (x"80",x"e0",x"c1",x"48"),
   329 => (x"bf",x"6e",x"7e",x"70"),
   330 => (x"87",x"c5",x"c0",x"02"),
   331 => (x"73",x"49",x"fe",x"4b"),
   332 => (x"48",x"a6",x"c8",x"0f"),
   333 => (x"fd",x"c3",x"78",x"c1"),
   334 => (x"87",x"db",x"e1",x"49"),
   335 => (x"99",x"c2",x"49",x"70"),
   336 => (x"87",x"e9",x"c0",x"02"),
   337 => (x"bf",x"d8",x"f5",x"c2"),
   338 => (x"87",x"c9",x"c0",x"02"),
   339 => (x"48",x"d8",x"f5",x"c2"),
   340 => (x"d3",x"c0",x"78",x"c0"),
   341 => (x"48",x"66",x"c4",x"87"),
   342 => (x"70",x"80",x"e0",x"c1"),
   343 => (x"02",x"bf",x"6e",x"7e"),
   344 => (x"4b",x"87",x"c5",x"c0"),
   345 => (x"0f",x"73",x"49",x"fd"),
   346 => (x"c1",x"48",x"a6",x"c8"),
   347 => (x"49",x"fa",x"c3",x"78"),
   348 => (x"70",x"87",x"e4",x"e0"),
   349 => (x"02",x"99",x"c2",x"49"),
   350 => (x"c2",x"87",x"ed",x"c0"),
   351 => (x"48",x"bf",x"d8",x"f5"),
   352 => (x"03",x"a8",x"b7",x"c7"),
   353 => (x"c2",x"87",x"c9",x"c0"),
   354 => (x"c7",x"48",x"d8",x"f5"),
   355 => (x"87",x"d3",x"c0",x"78"),
   356 => (x"c1",x"48",x"66",x"c4"),
   357 => (x"7e",x"70",x"80",x"e0"),
   358 => (x"c0",x"02",x"bf",x"6e"),
   359 => (x"fc",x"4b",x"87",x"c5"),
   360 => (x"c8",x"0f",x"73",x"49"),
   361 => (x"78",x"c1",x"48",x"a6"),
   362 => (x"f5",x"c2",x"7e",x"c0"),
   363 => (x"50",x"c0",x"48",x"d0"),
   364 => (x"c3",x"49",x"ee",x"cb"),
   365 => (x"a6",x"d4",x"87",x"c6"),
   366 => (x"d0",x"f5",x"c2",x"58"),
   367 => (x"c1",x"05",x"bf",x"97"),
   368 => (x"49",x"74",x"87",x"de"),
   369 => (x"05",x"99",x"f0",x"c3"),
   370 => (x"c1",x"87",x"cd",x"c0"),
   371 => (x"df",x"ff",x"49",x"da"),
   372 => (x"98",x"70",x"87",x"c5"),
   373 => (x"87",x"c8",x"c1",x"02"),
   374 => (x"bf",x"e8",x"7e",x"c1"),
   375 => (x"ff",x"c3",x"49",x"4b"),
   376 => (x"2b",x"b7",x"c8",x"99"),
   377 => (x"d9",x"c2",x"b3",x"71"),
   378 => (x"ff",x"49",x"bf",x"f8"),
   379 => (x"d0",x"87",x"e6",x"da"),
   380 => (x"d3",x"c2",x"49",x"66"),
   381 => (x"02",x"98",x"70",x"87"),
   382 => (x"c2",x"87",x"c6",x"c0"),
   383 => (x"c1",x"48",x"d0",x"f5"),
   384 => (x"d0",x"f5",x"c2",x"50"),
   385 => (x"c0",x"05",x"bf",x"97"),
   386 => (x"49",x"73",x"87",x"d6"),
   387 => (x"05",x"99",x"f0",x"c3"),
   388 => (x"c1",x"87",x"c5",x"ff"),
   389 => (x"dd",x"ff",x"49",x"da"),
   390 => (x"98",x"70",x"87",x"fd"),
   391 => (x"87",x"f8",x"fe",x"05"),
   392 => (x"e0",x"c0",x"02",x"6e"),
   393 => (x"48",x"a6",x"cc",x"87"),
   394 => (x"bf",x"d8",x"f5",x"c2"),
   395 => (x"49",x"66",x"cc",x"78"),
   396 => (x"66",x"c4",x"91",x"cc"),
   397 => (x"70",x"80",x"71",x"48"),
   398 => (x"02",x"bf",x"6e",x"7e"),
   399 => (x"4b",x"87",x"c6",x"c0"),
   400 => (x"73",x"49",x"66",x"cc"),
   401 => (x"02",x"66",x"c8",x"0f"),
   402 => (x"c2",x"87",x"c8",x"c0"),
   403 => (x"49",x"bf",x"d8",x"f5"),
   404 => (x"ec",x"87",x"e9",x"f1"),
   405 => (x"26",x"4d",x"26",x"8e"),
   406 => (x"26",x"4b",x"26",x"4c"),
   407 => (x"00",x"00",x"00",x"4f"),
   408 => (x"00",x"00",x"00",x"00"),
   409 => (x"14",x"11",x"12",x"58"),
   410 => (x"23",x"1c",x"1b",x"1d"),
   411 => (x"94",x"91",x"59",x"5a"),
   412 => (x"f4",x"eb",x"f2",x"f5"),
   413 => (x"00",x"00",x"00",x"00"),
   414 => (x"00",x"00",x"00",x"00"),
   415 => (x"ff",x"4a",x"71",x"1e"),
   416 => (x"72",x"49",x"bf",x"c8"),
   417 => (x"4f",x"26",x"48",x"a1"),
   418 => (x"bf",x"c8",x"ff",x"1e"),
   419 => (x"c0",x"c0",x"fe",x"89"),
   420 => (x"a9",x"c0",x"c0",x"c0"),
   421 => (x"c0",x"87",x"c4",x"01"),
   422 => (x"c1",x"87",x"c2",x"4a"),
   423 => (x"26",x"48",x"72",x"4a"),
   424 => (x"5b",x"5e",x"0e",x"4f"),
   425 => (x"71",x"0e",x"5d",x"5c"),
   426 => (x"4c",x"d4",x"ff",x"4b"),
   427 => (x"c0",x"48",x"66",x"d0"),
   428 => (x"ff",x"49",x"d6",x"78"),
   429 => (x"c3",x"87",x"dd",x"dd"),
   430 => (x"49",x"6c",x"7c",x"ff"),
   431 => (x"71",x"99",x"ff",x"c3"),
   432 => (x"f0",x"c3",x"49",x"4d"),
   433 => (x"a9",x"e0",x"c1",x"99"),
   434 => (x"c3",x"87",x"cb",x"05"),
   435 => (x"48",x"6c",x"7c",x"ff"),
   436 => (x"66",x"d0",x"98",x"c3"),
   437 => (x"ff",x"c3",x"78",x"08"),
   438 => (x"49",x"4a",x"6c",x"7c"),
   439 => (x"ff",x"c3",x"31",x"c8"),
   440 => (x"71",x"4a",x"6c",x"7c"),
   441 => (x"c8",x"49",x"72",x"b2"),
   442 => (x"7c",x"ff",x"c3",x"31"),
   443 => (x"b2",x"71",x"4a",x"6c"),
   444 => (x"31",x"c8",x"49",x"72"),
   445 => (x"6c",x"7c",x"ff",x"c3"),
   446 => (x"ff",x"b2",x"71",x"4a"),
   447 => (x"e0",x"c0",x"48",x"d0"),
   448 => (x"02",x"9b",x"73",x"78"),
   449 => (x"7b",x"72",x"87",x"c2"),
   450 => (x"4d",x"26",x"48",x"75"),
   451 => (x"4b",x"26",x"4c",x"26"),
   452 => (x"26",x"1e",x"4f",x"26"),
   453 => (x"5b",x"5e",x"0e",x"4f"),
   454 => (x"86",x"f8",x"0e",x"5c"),
   455 => (x"a6",x"c8",x"1e",x"76"),
   456 => (x"87",x"fd",x"fd",x"49"),
   457 => (x"4b",x"70",x"86",x"c4"),
   458 => (x"a8",x"c2",x"48",x"6e"),
   459 => (x"87",x"f0",x"c2",x"03"),
   460 => (x"f0",x"c3",x"4a",x"73"),
   461 => (x"aa",x"d0",x"c1",x"9a"),
   462 => (x"c1",x"87",x"c7",x"02"),
   463 => (x"c2",x"05",x"aa",x"e0"),
   464 => (x"49",x"73",x"87",x"de"),
   465 => (x"c3",x"02",x"99",x"c8"),
   466 => (x"87",x"c6",x"ff",x"87"),
   467 => (x"9c",x"c3",x"4c",x"73"),
   468 => (x"c1",x"05",x"ac",x"c2"),
   469 => (x"66",x"c4",x"87",x"c2"),
   470 => (x"71",x"31",x"c9",x"49"),
   471 => (x"4a",x"66",x"c4",x"1e"),
   472 => (x"f5",x"c2",x"92",x"d4"),
   473 => (x"81",x"72",x"49",x"dc"),
   474 => (x"87",x"e8",x"cd",x"fe"),
   475 => (x"da",x"ff",x"49",x"d8"),
   476 => (x"c0",x"c8",x"87",x"e2"),
   477 => (x"f4",x"e3",x"c2",x"1e"),
   478 => (x"da",x"e7",x"fd",x"49"),
   479 => (x"48",x"d0",x"ff",x"87"),
   480 => (x"c2",x"78",x"e0",x"c0"),
   481 => (x"cc",x"1e",x"f4",x"e3"),
   482 => (x"92",x"d4",x"4a",x"66"),
   483 => (x"49",x"dc",x"f5",x"c2"),
   484 => (x"cb",x"fe",x"81",x"72"),
   485 => (x"86",x"cc",x"87",x"ef"),
   486 => (x"c1",x"05",x"ac",x"c1"),
   487 => (x"66",x"c4",x"87",x"c2"),
   488 => (x"71",x"31",x"c9",x"49"),
   489 => (x"4a",x"66",x"c4",x"1e"),
   490 => (x"f5",x"c2",x"92",x"d4"),
   491 => (x"81",x"72",x"49",x"dc"),
   492 => (x"87",x"e0",x"cc",x"fe"),
   493 => (x"1e",x"f4",x"e3",x"c2"),
   494 => (x"d4",x"4a",x"66",x"c8"),
   495 => (x"dc",x"f5",x"c2",x"92"),
   496 => (x"fe",x"81",x"72",x"49"),
   497 => (x"d7",x"87",x"ef",x"c9"),
   498 => (x"c7",x"d9",x"ff",x"49"),
   499 => (x"1e",x"c0",x"c8",x"87"),
   500 => (x"49",x"f4",x"e3",x"c2"),
   501 => (x"87",x"dc",x"e5",x"fd"),
   502 => (x"d0",x"ff",x"86",x"cc"),
   503 => (x"78",x"e0",x"c0",x"48"),
   504 => (x"4c",x"26",x"8e",x"f8"),
   505 => (x"4f",x"26",x"4b",x"26"),
   506 => (x"5c",x"5b",x"5e",x"0e"),
   507 => (x"86",x"fc",x"0e",x"5d"),
   508 => (x"d4",x"ff",x"4d",x"71"),
   509 => (x"7e",x"66",x"d4",x"4c"),
   510 => (x"a8",x"b7",x"c3",x"48"),
   511 => (x"87",x"e2",x"c1",x"01"),
   512 => (x"66",x"c4",x"1e",x"75"),
   513 => (x"c2",x"93",x"d4",x"4b"),
   514 => (x"73",x"83",x"dc",x"f5"),
   515 => (x"e4",x"c3",x"fe",x"49"),
   516 => (x"49",x"a3",x"c8",x"87"),
   517 => (x"d0",x"ff",x"49",x"69"),
   518 => (x"78",x"e1",x"c8",x"48"),
   519 => (x"48",x"71",x"7c",x"dd"),
   520 => (x"70",x"98",x"ff",x"c3"),
   521 => (x"c8",x"4a",x"71",x"7c"),
   522 => (x"48",x"72",x"2a",x"b7"),
   523 => (x"70",x"98",x"ff",x"c3"),
   524 => (x"d0",x"4a",x"71",x"7c"),
   525 => (x"48",x"72",x"2a",x"b7"),
   526 => (x"70",x"98",x"ff",x"c3"),
   527 => (x"d8",x"48",x"71",x"7c"),
   528 => (x"7c",x"70",x"28",x"b7"),
   529 => (x"7c",x"7c",x"7c",x"c0"),
   530 => (x"7c",x"7c",x"7c",x"7c"),
   531 => (x"7c",x"7c",x"7c",x"7c"),
   532 => (x"48",x"d0",x"ff",x"7c"),
   533 => (x"c4",x"78",x"e0",x"c0"),
   534 => (x"49",x"dc",x"1e",x"66"),
   535 => (x"87",x"d9",x"d7",x"ff"),
   536 => (x"8e",x"fc",x"86",x"c8"),
   537 => (x"4c",x"26",x"4d",x"26"),
   538 => (x"4f",x"26",x"4b",x"26"),
   539 => (x"c0",x"1e",x"73",x"1e"),
   540 => (x"e2",x"c2",x"1e",x"4b"),
   541 => (x"fd",x"49",x"bf",x"e8"),
   542 => (x"86",x"c4",x"87",x"ee"),
   543 => (x"bf",x"ec",x"e2",x"c2"),
   544 => (x"c1",x"dc",x"fe",x"49"),
   545 => (x"05",x"98",x"70",x"87"),
   546 => (x"e2",x"c2",x"87",x"c4"),
   547 => (x"48",x"73",x"4b",x"d4"),
   548 => (x"4f",x"26",x"4b",x"26"),
   549 => (x"20",x"4d",x"4f",x"52"),
   550 => (x"64",x"61",x"6f",x"6c"),
   551 => (x"20",x"67",x"6e",x"69"),
   552 => (x"6c",x"69",x"61",x"66"),
   553 => (x"00",x"00",x"64",x"65"),
   554 => (x"00",x"00",x"28",x"b0"),
   555 => (x"00",x"00",x"28",x"bc"),
   556 => (x"20",x"43",x"42",x"42"),
   557 => (x"20",x"20",x"20",x"20"),
   558 => (x"00",x"44",x"48",x"56"),
   559 => (x"20",x"43",x"42",x"42"),
   560 => (x"20",x"20",x"20",x"20"),
   561 => (x"00",x"4d",x"4f",x"52"),
   562 => (x"00",x"00",x"1b",x"ab"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

