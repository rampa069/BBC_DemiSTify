library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c8f6c287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49c8f6c2",
    18 => x"48d0e3c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"d0e3c287",
    25 => x"cce3c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e8c187f7",
    29 => x"e3c287c6",
    30 => x"e3c24dd0",
    31 => x"ad744cd0",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"731e741e",
    65 => x"c11e721e",
    66 => x"87d0048b",
    67 => x"02114812",
    68 => x"c34c87ca",
    69 => x"749c98df",
    70 => x"87eb0288",
    71 => x"4b264a26",
    72 => x"4f264c26",
    73 => x"8148731e",
    74 => x"c502a973",
    75 => x"05531287",
    76 => x"4f2687f6",
    77 => x"711e731e",
    78 => x"4b66c84a",
    79 => x"718bc149",
    80 => x"87cf0299",
    81 => x"d4ff4812",
    82 => x"49737808",
    83 => x"99718bc1",
    84 => x"2687f105",
    85 => x"0e4f264b",
    86 => x"0e5c5b5e",
    87 => x"d4ff4a71",
    88 => x"4b66cc4c",
    89 => x"718bc149",
    90 => x"87ce0299",
    91 => x"6c7cffc3",
    92 => x"c1497352",
    93 => x"0599718b",
    94 => x"4c2687f2",
    95 => x"4f264b26",
    96 => x"ff1e731e",
    97 => x"ffc34bd4",
    98 => x"c34a6b7b",
    99 => x"496b7bff",
   100 => x"b17232c8",
   101 => x"6b7bffc3",
   102 => x"7131c84a",
   103 => x"7bffc3b2",
   104 => x"32c8496b",
   105 => x"4871b172",
   106 => x"4f264b26",
   107 => x"5c5b5e0e",
   108 => x"4d710e5d",
   109 => x"754cd4ff",
   110 => x"98ffc348",
   111 => x"e3c27c70",
   112 => x"c805bfd0",
   113 => x"4866d087",
   114 => x"a6d430c9",
   115 => x"4966d058",
   116 => x"487129d8",
   117 => x"7098ffc3",
   118 => x"4966d07c",
   119 => x"487129d0",
   120 => x"7098ffc3",
   121 => x"4966d07c",
   122 => x"487129c8",
   123 => x"7098ffc3",
   124 => x"4866d07c",
   125 => x"7098ffc3",
   126 => x"d049757c",
   127 => x"c3487129",
   128 => x"7c7098ff",
   129 => x"f0c94b6c",
   130 => x"ffc34aff",
   131 => x"87cf05ab",
   132 => x"6c7c7149",
   133 => x"028ac14b",
   134 => x"ab7187c5",
   135 => x"7387f202",
   136 => x"264d2648",
   137 => x"264b264c",
   138 => x"49c01e4f",
   139 => x"c348d4ff",
   140 => x"81c178ff",
   141 => x"a9b7c8c3",
   142 => x"2687f104",
   143 => x"5b5e0e4f",
   144 => x"c00e5d5c",
   145 => x"f7c1f0ff",
   146 => x"c0c0c14d",
   147 => x"4bc0c0c0",
   148 => x"c487d6ff",
   149 => x"c04cdff8",
   150 => x"fd49751e",
   151 => x"86c487ce",
   152 => x"c005a8c1",
   153 => x"d4ff87e5",
   154 => x"78ffc348",
   155 => x"e1c01e73",
   156 => x"49e9c1f0",
   157 => x"c487f5fc",
   158 => x"05987086",
   159 => x"d4ff87ca",
   160 => x"78ffc348",
   161 => x"87cb48c1",
   162 => x"c187defe",
   163 => x"c6ff058c",
   164 => x"2648c087",
   165 => x"264c264d",
   166 => x"0e4f264b",
   167 => x"0e5c5b5e",
   168 => x"c1f0ffc0",
   169 => x"d4ff4cc1",
   170 => x"78ffc348",
   171 => x"f749e0cb",
   172 => x"4bd387f5",
   173 => x"49741ec0",
   174 => x"c487f1fb",
   175 => x"05987086",
   176 => x"d4ff87ca",
   177 => x"78ffc348",
   178 => x"87cb48c1",
   179 => x"c187dafd",
   180 => x"dfff058b",
   181 => x"2648c087",
   182 => x"264b264c",
   183 => x"0000004f",
   184 => x"00444d43",
   185 => x"5c5b5e0e",
   186 => x"ffc30e5d",
   187 => x"4bd4ff4d",
   188 => x"c687f6fc",
   189 => x"e1c01eea",
   190 => x"49c8c1f0",
   191 => x"c487edfa",
   192 => x"02a8c186",
   193 => x"d2fe87c8",
   194 => x"c148c087",
   195 => x"eff987e8",
   196 => x"cf497087",
   197 => x"c699ffff",
   198 => x"c802a9ea",
   199 => x"87fbfd87",
   200 => x"d1c148c0",
   201 => x"c07b7587",
   202 => x"d0fc4cf1",
   203 => x"02987087",
   204 => x"c087ecc0",
   205 => x"f0ffc01e",
   206 => x"f949fac1",
   207 => x"86c487ee",
   208 => x"da059870",
   209 => x"6b7b7587",
   210 => x"757b7549",
   211 => x"757b757b",
   212 => x"99c0c17b",
   213 => x"c187c402",
   214 => x"c087db48",
   215 => x"c287d748",
   216 => x"87ca05ac",
   217 => x"f449c0ce",
   218 => x"48c087fd",
   219 => x"8cc187c8",
   220 => x"87f6fe05",
   221 => x"4d2648c0",
   222 => x"4b264c26",
   223 => x"00004f26",
   224 => x"43484453",
   225 => x"69616620",
   226 => x"000a216c",
   227 => x"5c5b5e0e",
   228 => x"d0ff0e5d",
   229 => x"d0e5c04d",
   230 => x"c24cc0c1",
   231 => x"c148d0e3",
   232 => x"49d8d078",
   233 => x"c787c0f4",
   234 => x"f97dc24b",
   235 => x"7dc387fb",
   236 => x"49741ec0",
   237 => x"c487f5f7",
   238 => x"05a8c186",
   239 => x"c24b87c1",
   240 => x"87cb05ab",
   241 => x"f349d0d0",
   242 => x"48c087dd",
   243 => x"c187f6c0",
   244 => x"d4ff058b",
   245 => x"87ccfc87",
   246 => x"58d4e3c2",
   247 => x"cd059870",
   248 => x"c01ec187",
   249 => x"d0c1f0ff",
   250 => x"87c0f749",
   251 => x"d4ff86c4",
   252 => x"78ffc348",
   253 => x"c287ccc5",
   254 => x"c258d8e3",
   255 => x"48d4ff7d",
   256 => x"c178ffc3",
   257 => x"264d2648",
   258 => x"264b264c",
   259 => x"0000004f",
   260 => x"52524549",
   261 => x"00000000",
   262 => x"00495053",
   263 => x"5c5b5e0e",
   264 => x"4d710e5d",
   265 => x"ff4cffc3",
   266 => x"7b744bd4",
   267 => x"c448d0ff",
   268 => x"7b7478c3",
   269 => x"ffc01e75",
   270 => x"49d8c1f0",
   271 => x"c487edf5",
   272 => x"02987086",
   273 => x"c8d287cb",
   274 => x"87dbf149",
   275 => x"eec048c1",
   276 => x"c37b7487",
   277 => x"c0c87bfe",
   278 => x"4966d41e",
   279 => x"c487d5f3",
   280 => x"747b7486",
   281 => x"d87b747b",
   282 => x"744ae0da",
   283 => x"c5056b7b",
   284 => x"058ac187",
   285 => x"7b7487f5",
   286 => x"c248d0ff",
   287 => x"2648c078",
   288 => x"264c264d",
   289 => x"004f264b",
   290 => x"74697257",
   291 => x"61662065",
   292 => x"64656c69",
   293 => x"5e0e000a",
   294 => x"0e5d5c5b",
   295 => x"4b7186fc",
   296 => x"c04cd4ff",
   297 => x"cdeec57e",
   298 => x"ffc34adf",
   299 => x"c3486c7c",
   300 => x"c005a8fe",
   301 => x"4d7487f8",
   302 => x"cc029b73",
   303 => x"1e66d487",
   304 => x"d2f24973",
   305 => x"d486c487",
   306 => x"48d0ff87",
   307 => x"d478d1c4",
   308 => x"ffc34a66",
   309 => x"058ac17d",
   310 => x"a6d887f8",
   311 => x"7cffc35a",
   312 => x"059b737c",
   313 => x"d0ff87c5",
   314 => x"c178d048",
   315 => x"8ac17e4a",
   316 => x"87f6fe05",
   317 => x"8efc486e",
   318 => x"4c264d26",
   319 => x"4f264b26",
   320 => x"711e731e",
   321 => x"ff4bc04a",
   322 => x"ffc348d4",
   323 => x"48d0ff78",
   324 => x"ff78c3c4",
   325 => x"ffc348d4",
   326 => x"c01e7278",
   327 => x"d1c1f0ff",
   328 => x"87c8f249",
   329 => x"987086c4",
   330 => x"c887d205",
   331 => x"66cc1ec0",
   332 => x"87e2fd49",
   333 => x"4b7086c4",
   334 => x"c248d0ff",
   335 => x"26487378",
   336 => x"0e4f264b",
   337 => x"5d5c5b5e",
   338 => x"c01ec00e",
   339 => x"c9c1f0ff",
   340 => x"87d8f149",
   341 => x"e3c21ed2",
   342 => x"f9fc49d8",
   343 => x"c086c887",
   344 => x"d284c14c",
   345 => x"f804acb7",
   346 => x"d8e3c287",
   347 => x"c349bf97",
   348 => x"c0c199c0",
   349 => x"e7c005a9",
   350 => x"dfe3c287",
   351 => x"d049bf97",
   352 => x"e0e3c231",
   353 => x"c84abf97",
   354 => x"c2b17232",
   355 => x"bf97e1e3",
   356 => x"4c71b14a",
   357 => x"ffffffcf",
   358 => x"ca84c19c",
   359 => x"87e7c134",
   360 => x"97e1e3c2",
   361 => x"31c149bf",
   362 => x"e3c299c6",
   363 => x"4abf97e2",
   364 => x"722ab7c7",
   365 => x"dde3c2b1",
   366 => x"4d4abf97",
   367 => x"e3c29dcf",
   368 => x"4abf97de",
   369 => x"32ca9ac3",
   370 => x"97dfe3c2",
   371 => x"33c24bbf",
   372 => x"e3c2b273",
   373 => x"4bbf97e0",
   374 => x"c69bc0c3",
   375 => x"b2732bb7",
   376 => x"48c181c2",
   377 => x"49703071",
   378 => x"307548c1",
   379 => x"4c724d70",
   380 => x"947184c1",
   381 => x"adb7c0c8",
   382 => x"c187cc06",
   383 => x"c82db734",
   384 => x"01adb7c0",
   385 => x"7487f4ff",
   386 => x"264d2648",
   387 => x"264b264c",
   388 => x"5b5e0e4f",
   389 => x"f80e5d5c",
   390 => x"c0ecc286",
   391 => x"c278c048",
   392 => x"c01ef8e3",
   393 => x"87d8fb49",
   394 => x"987086c4",
   395 => x"c087c505",
   396 => x"87c0c948",
   397 => x"7ec14dc0",
   398 => x"bfd8f7c0",
   399 => x"eee4c249",
   400 => x"4bc8714a",
   401 => x"7087dfea",
   402 => x"87c20598",
   403 => x"f7c07ec0",
   404 => x"c249bfd4",
   405 => x"714acae5",
   406 => x"c9ea4bc8",
   407 => x"05987087",
   408 => x"7ec087c2",
   409 => x"fdc0026e",
   410 => x"feeac287",
   411 => x"ebc24dbf",
   412 => x"7ebf9ff6",
   413 => x"ead6c548",
   414 => x"87c705a8",
   415 => x"bffeeac2",
   416 => x"6e87ce4d",
   417 => x"d5e9ca48",
   418 => x"87c502a8",
   419 => x"e3c748c0",
   420 => x"f8e3c287",
   421 => x"f949751e",
   422 => x"86c487e6",
   423 => x"c5059870",
   424 => x"c748c087",
   425 => x"f7c087ce",
   426 => x"c249bfd4",
   427 => x"714acae5",
   428 => x"f1e84bc8",
   429 => x"05987087",
   430 => x"ecc287c8",
   431 => x"78c148c0",
   432 => x"f7c087da",
   433 => x"c249bfd8",
   434 => x"714aeee4",
   435 => x"d5e84bc8",
   436 => x"02987087",
   437 => x"c087c5c0",
   438 => x"87d8c648",
   439 => x"97f6ebc2",
   440 => x"d5c149bf",
   441 => x"cdc005a9",
   442 => x"f7ebc287",
   443 => x"c249bf97",
   444 => x"c002a9ea",
   445 => x"48c087c5",
   446 => x"c287f9c5",
   447 => x"bf97f8e3",
   448 => x"e9c3487e",
   449 => x"cec002a8",
   450 => x"c3486e87",
   451 => x"c002a8eb",
   452 => x"48c087c5",
   453 => x"c287ddc5",
   454 => x"bf97c3e4",
   455 => x"c0059949",
   456 => x"e4c287cc",
   457 => x"49bf97c4",
   458 => x"c002a9c2",
   459 => x"48c087c5",
   460 => x"c287c1c5",
   461 => x"bf97c5e4",
   462 => x"fcebc248",
   463 => x"484c7058",
   464 => x"ecc288c1",
   465 => x"e4c258c0",
   466 => x"49bf97c6",
   467 => x"e4c28175",
   468 => x"4abf97c7",
   469 => x"a17232c8",
   470 => x"d0f0c27e",
   471 => x"c2786e48",
   472 => x"bf97c8e4",
   473 => x"58a6c848",
   474 => x"bfc0ecc2",
   475 => x"87cfc202",
   476 => x"bfd4f7c0",
   477 => x"cae5c249",
   478 => x"4bc8714a",
   479 => x"7087e7e5",
   480 => x"c5c00298",
   481 => x"c348c087",
   482 => x"ebc287ea",
   483 => x"c24cbff8",
   484 => x"c25ce4f0",
   485 => x"bf97dde4",
   486 => x"c231c849",
   487 => x"bf97dce4",
   488 => x"c249a14a",
   489 => x"bf97dee4",
   490 => x"7232d04a",
   491 => x"e4c249a1",
   492 => x"4abf97df",
   493 => x"a17232d8",
   494 => x"9166c449",
   495 => x"bfd0f0c2",
   496 => x"d8f0c281",
   497 => x"e5e4c259",
   498 => x"c84abf97",
   499 => x"e4e4c232",
   500 => x"a24bbf97",
   501 => x"e6e4c24a",
   502 => x"d04bbf97",
   503 => x"4aa27333",
   504 => x"97e7e4c2",
   505 => x"9bcf4bbf",
   506 => x"a27333d8",
   507 => x"dcf0c24a",
   508 => x"748ac25a",
   509 => x"dcf0c292",
   510 => x"78a17248",
   511 => x"c287c1c1",
   512 => x"bf97cae4",
   513 => x"c231c849",
   514 => x"bf97c9e4",
   515 => x"c549a14a",
   516 => x"81ffc731",
   517 => x"f0c229c9",
   518 => x"e4c259e4",
   519 => x"4abf97cf",
   520 => x"e4c232c8",
   521 => x"4bbf97ce",
   522 => x"66c44aa2",
   523 => x"c2826e92",
   524 => x"c25ae0f0",
   525 => x"c048d8f0",
   526 => x"d4f0c278",
   527 => x"78a17248",
   528 => x"48e4f0c2",
   529 => x"bfd8f0c2",
   530 => x"e8f0c278",
   531 => x"dcf0c248",
   532 => x"ecc278bf",
   533 => x"c002bfc0",
   534 => x"487487c9",
   535 => x"7e7030c4",
   536 => x"c287c9c0",
   537 => x"48bfe0f0",
   538 => x"7e7030c4",
   539 => x"48c4ecc2",
   540 => x"48c1786e",
   541 => x"4d268ef8",
   542 => x"4b264c26",
   543 => x"5e0e4f26",
   544 => x"0e5d5c5b",
   545 => x"ecc24a71",
   546 => x"cb02bfc0",
   547 => x"c74b7287",
   548 => x"c14d722b",
   549 => x"87c99dff",
   550 => x"2bc84b72",
   551 => x"ffc34d72",
   552 => x"d0f0c29d",
   553 => x"f7c083bf",
   554 => x"02abbfd0",
   555 => x"f7c087d9",
   556 => x"e3c25bd4",
   557 => x"49731ef8",
   558 => x"c487c5f1",
   559 => x"05987086",
   560 => x"48c087c5",
   561 => x"c287e6c0",
   562 => x"02bfc0ec",
   563 => x"497587d2",
   564 => x"e3c291c4",
   565 => x"4c6981f8",
   566 => x"ffffffcf",
   567 => x"87cb9cff",
   568 => x"91c24975",
   569 => x"81f8e3c2",
   570 => x"744c699f",
   571 => x"264d2648",
   572 => x"264b264c",
   573 => x"5b5e0e4f",
   574 => x"f40e5d5c",
   575 => x"59a6cc86",
   576 => x"c50566c8",
   577 => x"c348c087",
   578 => x"66c887c7",
   579 => x"7080c848",
   580 => x"78c0487e",
   581 => x"c70266dc",
   582 => x"9766dc87",
   583 => x"87c505bf",
   584 => x"ecc248c0",
   585 => x"c11ec087",
   586 => x"e9ca4949",
   587 => x"7086c487",
   588 => x"c0029c4c",
   589 => x"ecc287fc",
   590 => x"66dc4ac8",
   591 => x"cadeff49",
   592 => x"02987087",
   593 => x"7487ebc0",
   594 => x"4966dc4a",
   595 => x"deff4bcb",
   596 => x"987087ee",
   597 => x"c087db02",
   598 => x"029c741e",
   599 => x"4dc087c4",
   600 => x"4dc187c2",
   601 => x"edc94975",
   602 => x"7086c487",
   603 => x"ff059c4c",
   604 => x"9c7487c4",
   605 => x"87d7c102",
   606 => x"6e49a4dc",
   607 => x"da786948",
   608 => x"66c849a4",
   609 => x"c880c448",
   610 => x"699f58a6",
   611 => x"0866c448",
   612 => x"c0ecc278",
   613 => x"87d202bf",
   614 => x"9f49a4d4",
   615 => x"ffc04969",
   616 => x"487199ff",
   617 => x"7e7030d0",
   618 => x"7ec087c2",
   619 => x"66c4486e",
   620 => x"66c480bf",
   621 => x"66c87808",
   622 => x"c878c048",
   623 => x"81cc4966",
   624 => x"79bf66c4",
   625 => x"d04966c8",
   626 => x"c179c081",
   627 => x"c087c248",
   628 => x"268ef448",
   629 => x"264c264d",
   630 => x"0e4f264b",
   631 => x"5d5c5b5e",
   632 => x"d04c710e",
   633 => x"9c744d66",
   634 => x"87c2c102",
   635 => x"6949a4c8",
   636 => x"87fac002",
   637 => x"7585496c",
   638 => x"fcebc2b9",
   639 => x"baff4abf",
   640 => x"99719972",
   641 => x"87e4c002",
   642 => x"6b4ba4c4",
   643 => x"87eef949",
   644 => x"ebc27b70",
   645 => x"6c49bff8",
   646 => x"757c7181",
   647 => x"fcebc2b9",
   648 => x"baff4abf",
   649 => x"99719972",
   650 => x"87dcff05",
   651 => x"4d267c75",
   652 => x"4b264c26",
   653 => x"731e4f26",
   654 => x"9b4b711e",
   655 => x"c887c702",
   656 => x"056949a3",
   657 => x"48c087c5",
   658 => x"c287f6c0",
   659 => x"49bfd4f0",
   660 => x"6a4aa3c4",
   661 => x"c28ac24a",
   662 => x"92bff8eb",
   663 => x"c249a172",
   664 => x"4abffceb",
   665 => x"a1729a6b",
   666 => x"d4f7c049",
   667 => x"1e66c859",
   668 => x"87ccea71",
   669 => x"987086c4",
   670 => x"c087c405",
   671 => x"c187c248",
   672 => x"264b2648",
   673 => x"1e731e4f",
   674 => x"029b4b71",
   675 => x"a3c887c7",
   676 => x"c5056949",
   677 => x"c048c087",
   678 => x"f0c287f6",
   679 => x"c449bfd4",
   680 => x"4a6a4aa3",
   681 => x"ebc28ac2",
   682 => x"7292bff8",
   683 => x"ebc249a1",
   684 => x"6b4abffc",
   685 => x"49a1729a",
   686 => x"59d4f7c0",
   687 => x"711e66c8",
   688 => x"c487d9e5",
   689 => x"05987086",
   690 => x"48c087c4",
   691 => x"48c187c2",
   692 => x"4f264b26",
   693 => x"5c5b5e0e",
   694 => x"86fc0e5d",
   695 => x"66d44b71",
   696 => x"029b734d",
   697 => x"c887ccc1",
   698 => x"026949a3",
   699 => x"d087c4c1",
   700 => x"ebc24ca3",
   701 => x"ff49bffc",
   702 => x"994a6cb9",
   703 => x"a966d47e",
   704 => x"c087cd06",
   705 => x"a3cc7c7b",
   706 => x"49a3c44a",
   707 => x"87ca796a",
   708 => x"c0f84972",
   709 => x"4d66d499",
   710 => x"49758d71",
   711 => x"1e7129c9",
   712 => x"f6fa4973",
   713 => x"f8e3c287",
   714 => x"fc49731e",
   715 => x"86c887c8",
   716 => x"fc7c66d4",
   717 => x"264d268e",
   718 => x"264b264c",
   719 => x"1e731e4f",
   720 => x"029b4b71",
   721 => x"c287e4c0",
   722 => x"735be8f0",
   723 => x"c28ac24a",
   724 => x"49bff8eb",
   725 => x"d4f0c292",
   726 => x"807248bf",
   727 => x"58ecf0c2",
   728 => x"30c44871",
   729 => x"58c8ecc2",
   730 => x"c287edc0",
   731 => x"c248e4f0",
   732 => x"78bfd8f0",
   733 => x"48e8f0c2",
   734 => x"bfdcf0c2",
   735 => x"c0ecc278",
   736 => x"87c902bf",
   737 => x"bff8ebc2",
   738 => x"c731c449",
   739 => x"e0f0c287",
   740 => x"31c449bf",
   741 => x"59c8ecc2",
   742 => x"4f264b26",
   743 => x"5c5b5e0e",
   744 => x"c04a710e",
   745 => x"029a724b",
   746 => x"da87e0c0",
   747 => x"699f49a2",
   748 => x"c0ecc24b",
   749 => x"87cf02bf",
   750 => x"9f49a2d4",
   751 => x"c04c4969",
   752 => x"d09cffff",
   753 => x"c087c234",
   754 => x"73b3744c",
   755 => x"87edfd49",
   756 => x"4b264c26",
   757 => x"5e0e4f26",
   758 => x"0e5d5c5b",
   759 => x"a6c886f0",
   760 => x"ffffcf59",
   761 => x"c04cf8ff",
   762 => x"0266c47e",
   763 => x"e3c287d8",
   764 => x"78c048f4",
   765 => x"48ece3c2",
   766 => x"bfe8f0c2",
   767 => x"f0e3c278",
   768 => x"e4f0c248",
   769 => x"ecc278bf",
   770 => x"50c048d5",
   771 => x"bfc4ecc2",
   772 => x"f4e3c249",
   773 => x"aa714abf",
   774 => x"87cbc403",
   775 => x"99cf4972",
   776 => x"87e9c005",
   777 => x"48d0f7c0",
   778 => x"bfece3c2",
   779 => x"f8e3c278",
   780 => x"ece3c21e",
   781 => x"e3c249bf",
   782 => x"a1c148ec",
   783 => x"ffe27178",
   784 => x"c086c487",
   785 => x"c248ccf7",
   786 => x"cc78f8e3",
   787 => x"ccf7c087",
   788 => x"e0c048bf",
   789 => x"d0f7c080",
   790 => x"f4e3c258",
   791 => x"80c148bf",
   792 => x"58f8e3c2",
   793 => x"000dcc27",
   794 => x"bf97bf00",
   795 => x"c2029d4d",
   796 => x"e5c387e5",
   797 => x"dec202ad",
   798 => x"ccf7c087",
   799 => x"a3cb4bbf",
   800 => x"cf4c1149",
   801 => x"d2c105ac",
   802 => x"df497587",
   803 => x"cd89c199",
   804 => x"c8ecc291",
   805 => x"4aa3c181",
   806 => x"a3c35112",
   807 => x"c551124a",
   808 => x"51124aa3",
   809 => x"124aa3c7",
   810 => x"4aa3c951",
   811 => x"a3ce5112",
   812 => x"d051124a",
   813 => x"51124aa3",
   814 => x"124aa3d2",
   815 => x"4aa3d451",
   816 => x"a3d65112",
   817 => x"d851124a",
   818 => x"51124aa3",
   819 => x"124aa3dc",
   820 => x"4aa3de51",
   821 => x"7ec15112",
   822 => x"7487fcc0",
   823 => x"0599c849",
   824 => x"7487edc0",
   825 => x"0599d049",
   826 => x"e0c087d3",
   827 => x"ccc00266",
   828 => x"c0497387",
   829 => x"700f66e0",
   830 => x"d3c00298",
   831 => x"c0056e87",
   832 => x"ecc287c6",
   833 => x"50c048c8",
   834 => x"bfccf7c0",
   835 => x"87e9c248",
   836 => x"48d5ecc2",
   837 => x"c27e50c0",
   838 => x"49bfc4ec",
   839 => x"bff4e3c2",
   840 => x"04aa714a",
   841 => x"cf87f5fb",
   842 => x"f8ffffff",
   843 => x"e8f0c24c",
   844 => x"c8c005bf",
   845 => x"c0ecc287",
   846 => x"fac102bf",
   847 => x"f0e3c287",
   848 => x"f9ec49bf",
   849 => x"f4e3c287",
   850 => x"48a6c458",
   851 => x"bff0e3c2",
   852 => x"c0ecc278",
   853 => x"dbc002bf",
   854 => x"4966c487",
   855 => x"a9749974",
   856 => x"87c8c002",
   857 => x"c048a6c8",
   858 => x"87e7c078",
   859 => x"c148a6c8",
   860 => x"87dfc078",
   861 => x"cf4966c4",
   862 => x"a999f8ff",
   863 => x"87c8c002",
   864 => x"c048a6cc",
   865 => x"87c5c078",
   866 => x"c148a6cc",
   867 => x"48a6c878",
   868 => x"c87866cc",
   869 => x"dec00566",
   870 => x"4966c487",
   871 => x"ebc289c2",
   872 => x"c291bff8",
   873 => x"48bfd4f0",
   874 => x"e3c28071",
   875 => x"e3c258f0",
   876 => x"78c048f4",
   877 => x"c087d5f9",
   878 => x"ffffcf48",
   879 => x"f04cf8ff",
   880 => x"264d268e",
   881 => x"264b264c",
   882 => x"0000004f",
   883 => x"00000000",
   884 => x"ffffffff",
   885 => x"00000ddc",
   886 => x"00000de8",
   887 => x"33544146",
   888 => x"20202032",
   889 => x"00000000",
   890 => x"31544146",
   891 => x"20202036",
   892 => x"d4ff1e00",
   893 => x"78ffc348",
   894 => x"4f264868",
   895 => x"48d4ff1e",
   896 => x"ff78ffc3",
   897 => x"e1c048d0",
   898 => x"48d4ff78",
   899 => x"4f2678d4",
   900 => x"48d0ff1e",
   901 => x"2678e0c0",
   902 => x"d4ff1e4f",
   903 => x"99497087",
   904 => x"c087c602",
   905 => x"f105a9fb",
   906 => x"26487187",
   907 => x"5b5e0e4f",
   908 => x"4b710e5c",
   909 => x"f8fe4cc0",
   910 => x"99497087",
   911 => x"87f9c002",
   912 => x"02a9ecc0",
   913 => x"c087f2c0",
   914 => x"c002a9fb",
   915 => x"66cc87eb",
   916 => x"c703acb7",
   917 => x"0266d087",
   918 => x"537187c2",
   919 => x"c2029971",
   920 => x"fe84c187",
   921 => x"497087cb",
   922 => x"87cd0299",
   923 => x"02a9ecc0",
   924 => x"fbc087c7",
   925 => x"d5ff05a9",
   926 => x"0266d087",
   927 => x"97c087c3",
   928 => x"a9ecc07b",
   929 => x"7487c405",
   930 => x"7487c54a",
   931 => x"8a0ac04a",
   932 => x"4c264872",
   933 => x"4f264b26",
   934 => x"87d5fd1e",
   935 => x"c04a4970",
   936 => x"c904aaf0",
   937 => x"aaf9c087",
   938 => x"c087c301",
   939 => x"c1c18af0",
   940 => x"87c904aa",
   941 => x"01aadac1",
   942 => x"f7c087c3",
   943 => x"2648728a",
   944 => x"5b5e0e4f",
   945 => x"f80e5d5c",
   946 => x"c04c7186",
   947 => x"87ecfc7e",
   948 => x"fdc04bc0",
   949 => x"49bf97e0",
   950 => x"cf04a9c0",
   951 => x"87f9fc87",
   952 => x"fdc083c1",
   953 => x"49bf97e0",
   954 => x"87f106ab",
   955 => x"97e0fdc0",
   956 => x"87cf02bf",
   957 => x"7087fafb",
   958 => x"c6029949",
   959 => x"a9ecc087",
   960 => x"c087f105",
   961 => x"87e9fb4b",
   962 => x"e4fb4d70",
   963 => x"58a6c887",
   964 => x"7087defb",
   965 => x"c883c14a",
   966 => x"699749a4",
   967 => x"da05ad49",
   968 => x"49a4c987",
   969 => x"c4496997",
   970 => x"ce05a966",
   971 => x"49a4ca87",
   972 => x"aa496997",
   973 => x"c187c405",
   974 => x"c087d07e",
   975 => x"c602adec",
   976 => x"adfbc087",
   977 => x"c087c405",
   978 => x"6e7ec14b",
   979 => x"87f5fe02",
   980 => x"7387fdfa",
   981 => x"268ef848",
   982 => x"264c264d",
   983 => x"004f264b",
   984 => x"1e731e00",
   985 => x"c84bd4ff",
   986 => x"d0ff4a66",
   987 => x"78c5c848",
   988 => x"c148d4ff",
   989 => x"7b1178d4",
   990 => x"f9058ac1",
   991 => x"48d0ff87",
   992 => x"4b2678c4",
   993 => x"5e0e4f26",
   994 => x"0e5d5c5b",
   995 => x"7e7186f8",
   996 => x"f0c21e6e",
   997 => x"dce549f8",
   998 => x"7086c487",
   999 => x"e4c40298",
  1000 => x"e8ecc187",
  1001 => x"496e4cbf",
  1002 => x"c887d6fc",
  1003 => x"987058a6",
  1004 => x"c487c505",
  1005 => x"78c148a6",
  1006 => x"c548d0ff",
  1007 => x"48d4ff78",
  1008 => x"c478d5c1",
  1009 => x"89c14966",
  1010 => x"ecc131c6",
  1011 => x"4abf97e0",
  1012 => x"ffb07148",
  1013 => x"ff7808d4",
  1014 => x"78c448d0",
  1015 => x"97f4f0c2",
  1016 => x"99d049bf",
  1017 => x"c587dd02",
  1018 => x"48d4ff78",
  1019 => x"c078d6c1",
  1020 => x"48d4ff4a",
  1021 => x"c178ffc3",
  1022 => x"aae0c082",
  1023 => x"ff87f204",
  1024 => x"78c448d0",
  1025 => x"c348d4ff",
  1026 => x"d0ff78ff",
  1027 => x"ff78c548",
  1028 => x"d3c148d4",
  1029 => x"ff78c178",
  1030 => x"78c448d0",
  1031 => x"06acb7c0",
  1032 => x"c287cbc2",
  1033 => x"4bbfc0f1",
  1034 => x"737e748c",
  1035 => x"ddc1029b",
  1036 => x"4dc0c887",
  1037 => x"abb7c08b",
  1038 => x"c887c603",
  1039 => x"c04da3c0",
  1040 => x"f4f0c24b",
  1041 => x"d049bf97",
  1042 => x"87cf0299",
  1043 => x"f0c21ec0",
  1044 => x"e1e749f8",
  1045 => x"7086c487",
  1046 => x"c287d84c",
  1047 => x"c21ef8e3",
  1048 => x"e749f8f0",
  1049 => x"4c7087d0",
  1050 => x"e3c21e75",
  1051 => x"f0fb49f8",
  1052 => x"7486c887",
  1053 => x"87c5059c",
  1054 => x"cac148c0",
  1055 => x"c21ec187",
  1056 => x"e549f8f0",
  1057 => x"86c487d5",
  1058 => x"fe059b73",
  1059 => x"4c6e87e3",
  1060 => x"06acb7c0",
  1061 => x"f0c287d1",
  1062 => x"78c048f8",
  1063 => x"78c080d0",
  1064 => x"f1c280f4",
  1065 => x"c078bfc4",
  1066 => x"fd01acb7",
  1067 => x"d0ff87f5",
  1068 => x"ff78c548",
  1069 => x"d3c148d4",
  1070 => x"ff78c078",
  1071 => x"78c448d0",
  1072 => x"c2c048c1",
  1073 => x"f848c087",
  1074 => x"264d268e",
  1075 => x"264b264c",
  1076 => x"5b5e0e4f",
  1077 => x"fc0e5d5c",
  1078 => x"c04d7186",
  1079 => x"04ad4c4b",
  1080 => x"c087e8c0",
  1081 => x"741ec1fb",
  1082 => x"87c4029c",
  1083 => x"87c24ac0",
  1084 => x"49724ac1",
  1085 => x"c487dfeb",
  1086 => x"c17e7086",
  1087 => x"c2056e83",
  1088 => x"c14b7587",
  1089 => x"06ab7584",
  1090 => x"6e87d8ff",
  1091 => x"268efc48",
  1092 => x"264c264d",
  1093 => x"0e4f264b",
  1094 => x"0e5c5b5e",
  1095 => x"66cc4b71",
  1096 => x"4c87d802",
  1097 => x"028cf0c0",
  1098 => x"4a7487d8",
  1099 => x"d1028ac1",
  1100 => x"cd028a87",
  1101 => x"c9028a87",
  1102 => x"7387d987",
  1103 => x"87c6f949",
  1104 => x"1e7487d2",
  1105 => x"dac149c0",
  1106 => x"1e7487e2",
  1107 => x"dac14973",
  1108 => x"86c887da",
  1109 => x"4b264c26",
  1110 => x"5e0e4f26",
  1111 => x"0e5d5c5b",
  1112 => x"4c7186fc",
  1113 => x"c291de49",
  1114 => x"714de4f1",
  1115 => x"026d9785",
  1116 => x"c287dcc1",
  1117 => x"49bfd4f1",
  1118 => x"fd718174",
  1119 => x"7e7087d3",
  1120 => x"c0029848",
  1121 => x"f1c287f2",
  1122 => x"4a704bd8",
  1123 => x"fefe49cb",
  1124 => x"4b7487d2",
  1125 => x"ecc193cc",
  1126 => x"83c483ec",
  1127 => x"7bdcc7c1",
  1128 => x"c4c14974",
  1129 => x"7b7587da",
  1130 => x"97e4ecc1",
  1131 => x"c21e49bf",
  1132 => x"fd49d8f1",
  1133 => x"86c487e1",
  1134 => x"c4c14974",
  1135 => x"49c087c2",
  1136 => x"87ddc5c1",
  1137 => x"48f0f0c2",
  1138 => x"c04950c0",
  1139 => x"fc87cce2",
  1140 => x"264d268e",
  1141 => x"264b264c",
  1142 => x"0000004f",
  1143 => x"64616f4c",
  1144 => x"2e676e69",
  1145 => x"1e002e2e",
  1146 => x"4b711e73",
  1147 => x"d4f1c249",
  1148 => x"fb7181bf",
  1149 => x"4a7087db",
  1150 => x"87c4029a",
  1151 => x"87dce649",
  1152 => x"48d4f1c2",
  1153 => x"497378c0",
  1154 => x"2687fac1",
  1155 => x"1e4f264b",
  1156 => x"4b711e73",
  1157 => x"024aa3c4",
  1158 => x"c187d0c1",
  1159 => x"87dc028a",
  1160 => x"f2c0028a",
  1161 => x"c1058a87",
  1162 => x"f1c287d3",
  1163 => x"c102bfd4",
  1164 => x"c14887cb",
  1165 => x"d8f1c288",
  1166 => x"87c1c158",
  1167 => x"bfd4f1c2",
  1168 => x"c289c649",
  1169 => x"c059d8f1",
  1170 => x"c003a9b7",
  1171 => x"f1c287ef",
  1172 => x"78c048d4",
  1173 => x"c287e6c0",
  1174 => x"02bfd0f1",
  1175 => x"f1c287df",
  1176 => x"c148bfd4",
  1177 => x"d8f1c280",
  1178 => x"c287d258",
  1179 => x"02bfd0f1",
  1180 => x"f1c287cb",
  1181 => x"c648bfd4",
  1182 => x"d8f1c280",
  1183 => x"c4497358",
  1184 => x"264b2687",
  1185 => x"5b5e0e4f",
  1186 => x"f00e5d5c",
  1187 => x"59a6d086",
  1188 => x"4df8e3c2",
  1189 => x"f1c24cc0",
  1190 => x"78c148d0",
  1191 => x"c048a6c8",
  1192 => x"c27e7578",
  1193 => x"48bfd4f1",
  1194 => x"c106a8c0",
  1195 => x"a6c887c0",
  1196 => x"c27e755c",
  1197 => x"9848f8e3",
  1198 => x"87f2c002",
  1199 => x"c04d66c4",
  1200 => x"cc1ec1fb",
  1201 => x"87c40266",
  1202 => x"87c24cc0",
  1203 => x"49744cc1",
  1204 => x"c487c3e4",
  1205 => x"c17e7086",
  1206 => x"4866c885",
  1207 => x"a6cc80c1",
  1208 => x"d4f1c258",
  1209 => x"c503adbf",
  1210 => x"ff056e87",
  1211 => x"4d6e87d1",
  1212 => x"9d754cc0",
  1213 => x"87dcc302",
  1214 => x"1ec1fbc0",
  1215 => x"c70266cc",
  1216 => x"48a6c887",
  1217 => x"87c578c0",
  1218 => x"c148a6c8",
  1219 => x"4966c878",
  1220 => x"c487c3e3",
  1221 => x"487e7086",
  1222 => x"e4c20298",
  1223 => x"81cb4987",
  1224 => x"d0496997",
  1225 => x"d4c10299",
  1226 => x"cc497487",
  1227 => x"ececc191",
  1228 => x"e7c7c181",
  1229 => x"c381c879",
  1230 => x"497451ff",
  1231 => x"f1c291de",
  1232 => x"85714de4",
  1233 => x"7d97c1c2",
  1234 => x"c049a5c1",
  1235 => x"ecc251e0",
  1236 => x"02bf97c8",
  1237 => x"84c187d2",
  1238 => x"c24ba5c2",
  1239 => x"db4ac8ec",
  1240 => x"fff6fe49",
  1241 => x"87d9c187",
  1242 => x"c049a5cd",
  1243 => x"c284c151",
  1244 => x"4a6e4ba5",
  1245 => x"f6fe49cb",
  1246 => x"c4c187ea",
  1247 => x"cc497487",
  1248 => x"ececc191",
  1249 => x"dac5c181",
  1250 => x"c8ecc279",
  1251 => x"d802bf97",
  1252 => x"de497487",
  1253 => x"c284c191",
  1254 => x"714be4f1",
  1255 => x"c8ecc283",
  1256 => x"fe49dd4a",
  1257 => x"d887fdf5",
  1258 => x"de4b7487",
  1259 => x"e4f1c293",
  1260 => x"49a3cb83",
  1261 => x"84c151c0",
  1262 => x"cb4a6e73",
  1263 => x"e3f5fe49",
  1264 => x"4866c887",
  1265 => x"a6cc80c1",
  1266 => x"03acc758",
  1267 => x"6e87c5c0",
  1268 => x"87e4fc05",
  1269 => x"c003acc7",
  1270 => x"f1c287e4",
  1271 => x"78c048d0",
  1272 => x"91cc4974",
  1273 => x"81ececc1",
  1274 => x"79dac5c1",
  1275 => x"91de4974",
  1276 => x"81e4f1c2",
  1277 => x"84c151c0",
  1278 => x"ff04acc7",
  1279 => x"eec187dc",
  1280 => x"50c048c8",
  1281 => x"d1c180f7",
  1282 => x"d0c140f5",
  1283 => x"80c878e8",
  1284 => x"78cfc8c1",
  1285 => x"c04966cc",
  1286 => x"f087e5fa",
  1287 => x"264d268e",
  1288 => x"264b264c",
  1289 => x"0000004f",
  1290 => x"61422080",
  1291 => x"1e006b63",
  1292 => x"4b711e73",
  1293 => x"c191cc49",
  1294 => x"c881ecec",
  1295 => x"ecc14aa1",
  1296 => x"501248e0",
  1297 => x"c04aa1c9",
  1298 => x"1248e0fd",
  1299 => x"c181ca50",
  1300 => x"1148e4ec",
  1301 => x"e4ecc150",
  1302 => x"1e49bf97",
  1303 => x"f6f249c0",
  1304 => x"f8497387",
  1305 => x"8efc87df",
  1306 => x"4f264b26",
  1307 => x"c049c01e",
  1308 => x"2687eefa",
  1309 => x"4a711e4f",
  1310 => x"c191cc49",
  1311 => x"c881ecec",
  1312 => x"f0f0c281",
  1313 => x"c0501148",
  1314 => x"fe49a2f0",
  1315 => x"c087fdef",
  1316 => x"87c7d749",
  1317 => x"ff1e4f26",
  1318 => x"ffc34ad4",
  1319 => x"48d0ff7a",
  1320 => x"de78e1c0",
  1321 => x"487a717a",
  1322 => x"7028b7c8",
  1323 => x"d048717a",
  1324 => x"7a7028b7",
  1325 => x"b7d84871",
  1326 => x"ff7a7028",
  1327 => x"e0c048d0",
  1328 => x"0e4f2678",
  1329 => x"5d5c5b5e",
  1330 => x"7186f40e",
  1331 => x"91cc494d",
  1332 => x"81ececc1",
  1333 => x"ca4aa1c8",
  1334 => x"a6c47ea1",
  1335 => x"ecf0c248",
  1336 => x"976e78bf",
  1337 => x"66c44bbf",
  1338 => x"122c734c",
  1339 => x"58a6cc48",
  1340 => x"84c19c70",
  1341 => x"699781c9",
  1342 => x"04acb749",
  1343 => x"4cc087c2",
  1344 => x"4abf976e",
  1345 => x"724966c8",
  1346 => x"c4b9ff31",
  1347 => x"48749966",
  1348 => x"4a703072",
  1349 => x"f0f0c2b1",
  1350 => x"f9fd7159",
  1351 => x"c21ec787",
  1352 => x"1ebfccf1",
  1353 => x"1eececc1",
  1354 => x"97f0f0c2",
  1355 => x"f4c149bf",
  1356 => x"c0497587",
  1357 => x"e887c9f6",
  1358 => x"264d268e",
  1359 => x"264b264c",
  1360 => x"1e731e4f",
  1361 => x"fd494b71",
  1362 => x"497387f9",
  1363 => x"2687f4fd",
  1364 => x"1e4f264b",
  1365 => x"4b711e73",
  1366 => x"024aa3c2",
  1367 => x"8ac187d6",
  1368 => x"87e2c005",
  1369 => x"bfccf1c2",
  1370 => x"4887db02",
  1371 => x"f1c288c1",
  1372 => x"87d258d0",
  1373 => x"bfd0f1c2",
  1374 => x"c287cb02",
  1375 => x"48bfccf1",
  1376 => x"f1c280c1",
  1377 => x"1ec758d0",
  1378 => x"bfccf1c2",
  1379 => x"ececc11e",
  1380 => x"f0f0c21e",
  1381 => x"cc49bf97",
  1382 => x"c0497387",
  1383 => x"f487e1f4",
  1384 => x"264b268e",
  1385 => x"5b5e0e4f",
  1386 => x"ff0e5d5c",
  1387 => x"e4c086cc",
  1388 => x"a6cc59a6",
  1389 => x"c478c048",
  1390 => x"c478c080",
  1391 => x"66c8c180",
  1392 => x"c180c478",
  1393 => x"c180c478",
  1394 => x"d0f1c278",
  1395 => x"e078c148",
  1396 => x"c4e187ea",
  1397 => x"87d9e087",
  1398 => x"fbc04c70",
  1399 => x"f3c102ac",
  1400 => x"66e0c087",
  1401 => x"87e8c105",
  1402 => x"4a66c4c1",
  1403 => x"7e6a82c4",
  1404 => x"48fce8c1",
  1405 => x"4120496e",
  1406 => x"51104120",
  1407 => x"4866c4c1",
  1408 => x"78efd0c1",
  1409 => x"81c7496a",
  1410 => x"c4c15174",
  1411 => x"81c84966",
  1412 => x"a6d851c1",
  1413 => x"c178c248",
  1414 => x"c94966c4",
  1415 => x"c151c081",
  1416 => x"ca4966c4",
  1417 => x"c151c081",
  1418 => x"6a1ed81e",
  1419 => x"ff81c849",
  1420 => x"c887fadf",
  1421 => x"66c8c186",
  1422 => x"01a8c048",
  1423 => x"a6d087c7",
  1424 => x"cf78c148",
  1425 => x"66c8c187",
  1426 => x"d888c148",
  1427 => x"87c458a6",
  1428 => x"87c5dfff",
  1429 => x"cd029c74",
  1430 => x"66d087da",
  1431 => x"66ccc148",
  1432 => x"cfcd03a8",
  1433 => x"48a6c887",
  1434 => x"ff7e78c0",
  1435 => x"7087c2de",
  1436 => x"acd0c14c",
  1437 => x"87e7c205",
  1438 => x"6e48a6c4",
  1439 => x"87d8e078",
  1440 => x"cc487e70",
  1441 => x"c506a866",
  1442 => x"48a6cc87",
  1443 => x"ddff786e",
  1444 => x"4c7087df",
  1445 => x"05acecc0",
  1446 => x"d087eec1",
  1447 => x"91cc4966",
  1448 => x"8166c4c1",
  1449 => x"6a4aa1c4",
  1450 => x"4aa1c84d",
  1451 => x"d1c1526e",
  1452 => x"dcff79f5",
  1453 => x"4c7087fb",
  1454 => x"87d9029c",
  1455 => x"02acfbc0",
  1456 => x"557487d3",
  1457 => x"87e9dcff",
  1458 => x"029c4c70",
  1459 => x"fbc087c7",
  1460 => x"edff05ac",
  1461 => x"55e0c087",
  1462 => x"c055c1c2",
  1463 => x"e0c07d97",
  1464 => x"66c44866",
  1465 => x"87db05a8",
  1466 => x"d44866d0",
  1467 => x"ca04a866",
  1468 => x"4866d087",
  1469 => x"a6d480c1",
  1470 => x"d487c858",
  1471 => x"88c14866",
  1472 => x"ff58a6d8",
  1473 => x"7087eadb",
  1474 => x"acd0c14c",
  1475 => x"dc87c905",
  1476 => x"80c14866",
  1477 => x"58a6e0c0",
  1478 => x"02acd0c1",
  1479 => x"6e87d9fd",
  1480 => x"66e0c048",
  1481 => x"ebc905a8",
  1482 => x"a6e4c087",
  1483 => x"7478c048",
  1484 => x"88fbc048",
  1485 => x"7058a6c8",
  1486 => x"ddc90298",
  1487 => x"88cb4887",
  1488 => x"7058a6c8",
  1489 => x"cfc10298",
  1490 => x"88c94887",
  1491 => x"7058a6c8",
  1492 => x"ffc30298",
  1493 => x"88c44887",
  1494 => x"7058a6c8",
  1495 => x"87cf0298",
  1496 => x"c888c148",
  1497 => x"987058a6",
  1498 => x"87e8c302",
  1499 => x"c887dcc8",
  1500 => x"f0c048a6",
  1501 => x"f8d9ff78",
  1502 => x"c04c7087",
  1503 => x"c002acec",
  1504 => x"a6cc87c3",
  1505 => x"acecc05c",
  1506 => x"ff87cd02",
  1507 => x"7087e2d9",
  1508 => x"acecc04c",
  1509 => x"87f3ff05",
  1510 => x"02acecc0",
  1511 => x"ff87c4c0",
  1512 => x"c087ced9",
  1513 => x"d81eca1e",
  1514 => x"91cc4966",
  1515 => x"4866ccc1",
  1516 => x"a6cc8071",
  1517 => x"4866c858",
  1518 => x"a6d080c4",
  1519 => x"bf66cc58",
  1520 => x"e8d9ff49",
  1521 => x"de1ec187",
  1522 => x"bf66d41e",
  1523 => x"dcd9ff49",
  1524 => x"7086d087",
  1525 => x"08c04849",
  1526 => x"a6ecc088",
  1527 => x"06a8c058",
  1528 => x"c087eec0",
  1529 => x"dd4866e8",
  1530 => x"e4c003a8",
  1531 => x"bf66c487",
  1532 => x"66e8c049",
  1533 => x"51e0c081",
  1534 => x"4966e8c0",
  1535 => x"66c481c1",
  1536 => x"c1c281bf",
  1537 => x"66e8c051",
  1538 => x"c481c249",
  1539 => x"c081bf66",
  1540 => x"c1486e51",
  1541 => x"6e78efd0",
  1542 => x"d881c849",
  1543 => x"496e5166",
  1544 => x"66dc81c9",
  1545 => x"ca496e51",
  1546 => x"5166c881",
  1547 => x"c14866d8",
  1548 => x"58a6dc80",
  1549 => x"d44866d0",
  1550 => x"c004a866",
  1551 => x"66d087cb",
  1552 => x"d480c148",
  1553 => x"d1c558a6",
  1554 => x"4866d487",
  1555 => x"a6d888c1",
  1556 => x"87c6c558",
  1557 => x"87c0d9ff",
  1558 => x"58a6ecc0",
  1559 => x"87f8d8ff",
  1560 => x"58a6f0c0",
  1561 => x"05a8ecc0",
  1562 => x"a687c9c0",
  1563 => x"66e8c048",
  1564 => x"87c4c078",
  1565 => x"87f9d5ff",
  1566 => x"cc4966d0",
  1567 => x"66c4c191",
  1568 => x"c8807148",
  1569 => x"66c458a6",
  1570 => x"c482c84a",
  1571 => x"81ca4966",
  1572 => x"5166e8c0",
  1573 => x"4966ecc0",
  1574 => x"e8c081c1",
  1575 => x"48c18966",
  1576 => x"49703071",
  1577 => x"977189c1",
  1578 => x"ecf0c27a",
  1579 => x"e8c049bf",
  1580 => x"6a972966",
  1581 => x"9871484a",
  1582 => x"58a6f4c0",
  1583 => x"c44866c4",
  1584 => x"58a6cc80",
  1585 => x"4dbf66c8",
  1586 => x"4866e0c0",
  1587 => x"c002a86e",
  1588 => x"7ec087c5",
  1589 => x"c187c2c0",
  1590 => x"c01e6e7e",
  1591 => x"49751ee0",
  1592 => x"87c9d5ff",
  1593 => x"4c7086c8",
  1594 => x"06acb7c0",
  1595 => x"7487d4c1",
  1596 => x"bf66c885",
  1597 => x"81e0c049",
  1598 => x"c14b8975",
  1599 => x"714ac8e9",
  1600 => x"87e0e0fe",
  1601 => x"7e7585c2",
  1602 => x"4866e4c0",
  1603 => x"e8c080c1",
  1604 => x"f0c058a6",
  1605 => x"81c14966",
  1606 => x"c002a970",
  1607 => x"4dc087c5",
  1608 => x"c187c2c0",
  1609 => x"cc1e754d",
  1610 => x"c049bf66",
  1611 => x"66c481e0",
  1612 => x"c81e7189",
  1613 => x"d3ff4966",
  1614 => x"86c887f3",
  1615 => x"01a8b7c0",
  1616 => x"c087c5ff",
  1617 => x"c00266e4",
  1618 => x"66c487d3",
  1619 => x"c081c949",
  1620 => x"c45166e4",
  1621 => x"d3c14866",
  1622 => x"cec078c3",
  1623 => x"4966c487",
  1624 => x"51c281c9",
  1625 => x"c14866c4",
  1626 => x"d078c1d5",
  1627 => x"66d44866",
  1628 => x"cbc004a8",
  1629 => x"4866d087",
  1630 => x"a6d480c1",
  1631 => x"87dac058",
  1632 => x"c14866d4",
  1633 => x"58a6d888",
  1634 => x"ff87cfc0",
  1635 => x"7087cad2",
  1636 => x"87c6c04c",
  1637 => x"87c1d2ff",
  1638 => x"66dc4c70",
  1639 => x"c080c148",
  1640 => x"7458a6e0",
  1641 => x"cbc0029c",
  1642 => x"4866d087",
  1643 => x"a866ccc1",
  1644 => x"87f1f204",
  1645 => x"c74866d0",
  1646 => x"e1c003a8",
  1647 => x"4c66d087",
  1648 => x"48d0f1c2",
  1649 => x"497478c0",
  1650 => x"c4c191cc",
  1651 => x"a1c48166",
  1652 => x"c04a6a4a",
  1653 => x"84c17952",
  1654 => x"ff04acc7",
  1655 => x"e0c087e2",
  1656 => x"e2c00266",
  1657 => x"66c4c187",
  1658 => x"81d4c149",
  1659 => x"4a66c4c1",
  1660 => x"c082dcc1",
  1661 => x"f5d1c152",
  1662 => x"66c4c179",
  1663 => x"81d8c149",
  1664 => x"79cce9c1",
  1665 => x"c187d6c0",
  1666 => x"c14966c4",
  1667 => x"c4c181d4",
  1668 => x"d8c14a66",
  1669 => x"d4e9c182",
  1670 => x"ecd1c17a",
  1671 => x"66c4c179",
  1672 => x"81e0c149",
  1673 => x"79d3d5c1",
  1674 => x"87e4cfff",
  1675 => x"ff4866cc",
  1676 => x"4d268ecc",
  1677 => x"4b264c26",
  1678 => x"00004f26",
  1679 => x"64616f4c",
  1680 => x"202e2a20",
  1681 => x"00000000",
  1682 => x"0000203a",
  1683 => x"61422080",
  1684 => x"00006b63",
  1685 => x"78452080",
  1686 => x"1e007469",
  1687 => x"f1c21ec7",
  1688 => x"c11ebfcc",
  1689 => x"c21eecec",
  1690 => x"bf97f0f0",
  1691 => x"87f5ec49",
  1692 => x"49ececc1",
  1693 => x"87d6e2c0",
  1694 => x"4f268ef4",
  1695 => x"c81e731e",
  1696 => x"eec187c3",
  1697 => x"ecc148c4",
  1698 => x"e8fe78cc",
  1699 => x"e1c049a0",
  1700 => x"49c787fc",
  1701 => x"87e8e0c0",
  1702 => x"e2c049c1",
  1703 => x"d4ff87c3",
  1704 => x"78ffc348",
  1705 => x"48d8f1c2",
  1706 => x"e3fe50c0",
  1707 => x"987087de",
  1708 => x"fe87cd02",
  1709 => x"7087daed",
  1710 => x"87c40298",
  1711 => x"87c24ac1",
  1712 => x"9a724ac0",
  1713 => x"c187c802",
  1714 => x"fe49d8ec",
  1715 => x"c287d8d7",
  1716 => x"c048ccf1",
  1717 => x"f0f0c278",
  1718 => x"4950c048",
  1719 => x"c087fcfd",
  1720 => x"7087cdf6",
  1721 => x"cb029b4b",
  1722 => x"c8eec187",
  1723 => x"df49c75b",
  1724 => x"87c687ce",
  1725 => x"e0c049c0",
  1726 => x"c2c387e7",
  1727 => x"c8e2c087",
  1728 => x"d4f0c087",
  1729 => x"87f5ff87",
  1730 => x"4f264b26",
  1731 => x"746f6f42",
  1732 => x"2e676e69",
  1733 => x"00002e2e",
  1734 => x"4f204453",
  1735 => x"0000004b",
  1736 => x"00000000",
  1737 => x"00000000",
  1738 => x"00000001",
  1739 => x"0000115a",
  1740 => x"00002c64",
  1741 => x"00000000",
  1742 => x"0000115a",
  1743 => x"00002c82",
  1744 => x"00000000",
  1745 => x"0000115a",
  1746 => x"00002ca0",
  1747 => x"00000000",
  1748 => x"0000115a",
  1749 => x"00002cbe",
  1750 => x"00000000",
  1751 => x"0000115a",
  1752 => x"00002cdc",
  1753 => x"00000000",
  1754 => x"0000115a",
  1755 => x"00002cfa",
  1756 => x"00000000",
  1757 => x"0000115a",
  1758 => x"00002d18",
  1759 => x"00000000",
  1760 => x"00001475",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"0000120f",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"db86fc1e",
  1767 => x"fc7e7087",
  1768 => x"1e4f268e",
  1769 => x"c048f0fe",
  1770 => x"7909cd78",
  1771 => x"1e4f2609",
  1772 => x"49d8eec1",
  1773 => x"4f2687ed",
  1774 => x"bff0fe1e",
  1775 => x"1e4f2648",
  1776 => x"c148f0fe",
  1777 => x"1e4f2678",
  1778 => x"c048f0fe",
  1779 => x"1e4f2678",
  1780 => x"52c04a71",
  1781 => x"0e4f2651",
  1782 => x"5d5c5b5e",
  1783 => x"7186f40e",
  1784 => x"7e6d974d",
  1785 => x"974ca5c1",
  1786 => x"a6c8486c",
  1787 => x"c4486e58",
  1788 => x"c505a866",
  1789 => x"c048ff87",
  1790 => x"caff87e6",
  1791 => x"49a5c287",
  1792 => x"714b6c97",
  1793 => x"6b974ba3",
  1794 => x"7e6c974b",
  1795 => x"80c1486e",
  1796 => x"c758a6c8",
  1797 => x"58a6cc98",
  1798 => x"fe7c9770",
  1799 => x"487387e1",
  1800 => x"4d268ef4",
  1801 => x"4b264c26",
  1802 => x"5e0e4f26",
  1803 => x"f40e5c5b",
  1804 => x"d84c7186",
  1805 => x"ffc34a66",
  1806 => x"4ba4c29a",
  1807 => x"73496c97",
  1808 => x"517249a1",
  1809 => x"6e7e6c97",
  1810 => x"c880c148",
  1811 => x"98c758a6",
  1812 => x"7058a6cc",
  1813 => x"268ef454",
  1814 => x"264b264c",
  1815 => x"86fc1e4f",
  1816 => x"e087e4fd",
  1817 => x"c0494abf",
  1818 => x"0299c0e0",
  1819 => x"1e7287cb",
  1820 => x"49f8f4c2",
  1821 => x"c487f3fe",
  1822 => x"87fcfc86",
  1823 => x"fefc7e70",
  1824 => x"268efc87",
  1825 => x"f4c21e4f",
  1826 => x"c2fd49f8",
  1827 => x"ddf1c187",
  1828 => x"87cffc49",
  1829 => x"2687edc3",
  1830 => x"5b5e0e4f",
  1831 => x"fc0e5d5c",
  1832 => x"ff7e7186",
  1833 => x"f4c24dd4",
  1834 => x"eafc49f8",
  1835 => x"c04b7087",
  1836 => x"c204abb7",
  1837 => x"f0c387f8",
  1838 => x"87c905ab",
  1839 => x"48fcf5c1",
  1840 => x"d9c278c1",
  1841 => x"abe0c387",
  1842 => x"c187c905",
  1843 => x"c148c0f6",
  1844 => x"87cac278",
  1845 => x"bfc0f6c1",
  1846 => x"c287c602",
  1847 => x"c24ca3c0",
  1848 => x"c14c7387",
  1849 => x"02bffcf5",
  1850 => x"7487e0c0",
  1851 => x"29b7c449",
  1852 => x"d8f7c191",
  1853 => x"cf4a7481",
  1854 => x"c192c29a",
  1855 => x"70307248",
  1856 => x"72baff4a",
  1857 => x"70986948",
  1858 => x"7487db79",
  1859 => x"29b7c449",
  1860 => x"d8f7c191",
  1861 => x"cf4a7481",
  1862 => x"c392c29a",
  1863 => x"70307248",
  1864 => x"b069484a",
  1865 => x"056e7970",
  1866 => x"ff87e7c0",
  1867 => x"e1c848d0",
  1868 => x"c17dc578",
  1869 => x"02bfc0f6",
  1870 => x"e0c387c3",
  1871 => x"fcf5c17d",
  1872 => x"87c302bf",
  1873 => x"737df0c3",
  1874 => x"48d0ff7d",
  1875 => x"c078e1c8",
  1876 => x"f6c178e0",
  1877 => x"78c048c0",
  1878 => x"48fcf5c1",
  1879 => x"f4c278c0",
  1880 => x"f2f949f8",
  1881 => x"c04b7087",
  1882 => x"fd03abb7",
  1883 => x"48c087c8",
  1884 => x"4d268efc",
  1885 => x"4b264c26",
  1886 => x"00004f26",
  1887 => x"00000000",
  1888 => x"00000000",
  1889 => x"724ac01e",
  1890 => x"c191c449",
  1891 => x"c081d8f7",
  1892 => x"d082c179",
  1893 => x"ee04aab7",
  1894 => x"0e4f2687",
  1895 => x"5d5c5b5e",
  1896 => x"f84d710e",
  1897 => x"4a7587e1",
  1898 => x"922ab7c4",
  1899 => x"82d8f7c1",
  1900 => x"9ccf4c75",
  1901 => x"496a94c2",
  1902 => x"c32b744b",
  1903 => x"7448c29b",
  1904 => x"ff4c7030",
  1905 => x"714874bc",
  1906 => x"f77a7098",
  1907 => x"487387f1",
  1908 => x"4c264d26",
  1909 => x"4f264b26",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"00000000",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"00000000",
  1926 => x"48d0ff1e",
  1927 => x"7178e1c8",
  1928 => x"08d4ff48",
  1929 => x"1e4f2678",
  1930 => x"c848d0ff",
  1931 => x"487178e1",
  1932 => x"7808d4ff",
  1933 => x"ff4866c4",
  1934 => x"267808d4",
  1935 => x"4a711e4f",
  1936 => x"1e4966c4",
  1937 => x"deff4972",
  1938 => x"48d0ff87",
  1939 => x"fc78e0c0",
  1940 => x"1e4f268e",
  1941 => x"4b711e73",
  1942 => x"1e4966c8",
  1943 => x"e0c14a73",
  1944 => x"d8ff49a2",
  1945 => x"268efc87",
  1946 => x"1e4f264b",
  1947 => x"c848d0ff",
  1948 => x"487178c9",
  1949 => x"7808d4ff",
  1950 => x"711e4f26",
  1951 => x"87eb494a",
  1952 => x"c848d0ff",
  1953 => x"1e4f2678",
  1954 => x"4b711e73",
  1955 => x"bfd0f5c2",
  1956 => x"c287c302",
  1957 => x"d0ff87eb",
  1958 => x"78c9c848",
  1959 => x"e0c04873",
  1960 => x"08d4ffb0",
  1961 => x"c4f5c278",
  1962 => x"c878c048",
  1963 => x"87c50266",
  1964 => x"c249ffc3",
  1965 => x"c249c087",
  1966 => x"cc59ccf5",
  1967 => x"87c60266",
  1968 => x"4ad5d5c5",
  1969 => x"ffcf87c4",
  1970 => x"f5c24aff",
  1971 => x"f5c25ad0",
  1972 => x"78c148d0",
  1973 => x"4f264b26",
  1974 => x"5c5b5e0e",
  1975 => x"4d710e5d",
  1976 => x"bfccf5c2",
  1977 => x"029d754b",
  1978 => x"c84987cb",
  1979 => x"c0fac191",
  1980 => x"c482714a",
  1981 => x"c0fec187",
  1982 => x"124cc04a",
  1983 => x"c2997349",
  1984 => x"48bfc8f5",
  1985 => x"d4ffb871",
  1986 => x"b7c17808",
  1987 => x"b7c8842b",
  1988 => x"87e704ac",
  1989 => x"bfc4f5c2",
  1990 => x"c280c848",
  1991 => x"2658c8f5",
  1992 => x"264c264d",
  1993 => x"1e4f264b",
  1994 => x"4b711e73",
  1995 => x"029a4a13",
  1996 => x"497287cb",
  1997 => x"1387e1fe",
  1998 => x"f5059a4a",
  1999 => x"264b2687",
  2000 => x"f5c21e4f",
  2001 => x"c249bfc4",
  2002 => x"c148c4f5",
  2003 => x"c0c478a1",
  2004 => x"db03a9b7",
  2005 => x"48d4ff87",
  2006 => x"bfc8f5c2",
  2007 => x"c4f5c278",
  2008 => x"f5c249bf",
  2009 => x"a1c148c4",
  2010 => x"b7c0c478",
  2011 => x"87e504a9",
  2012 => x"c848d0ff",
  2013 => x"d0f5c278",
  2014 => x"2678c048",
  2015 => x"0000004f",
  2016 => x"00000000",
  2017 => x"00000000",
  2018 => x"5f000000",
  2019 => x"0000005f",
  2020 => x"00030300",
  2021 => x"00000303",
  2022 => x"147f7f14",
  2023 => x"00147f7f",
  2024 => x"6b2e2400",
  2025 => x"00123a6b",
  2026 => x"18366a4c",
  2027 => x"0032566c",
  2028 => x"594f7e30",
  2029 => x"40683a77",
  2030 => x"07040000",
  2031 => x"00000003",
  2032 => x"3e1c0000",
  2033 => x"00004163",
  2034 => x"63410000",
  2035 => x"00001c3e",
  2036 => x"1c3e2a08",
  2037 => x"082a3e1c",
  2038 => x"3e080800",
  2039 => x"0008083e",
  2040 => x"e0800000",
  2041 => x"00000060",
  2042 => x"08080800",
  2043 => x"00080808",
  2044 => x"60000000",
  2045 => x"00000060",
  2046 => x"18306040",
  2047 => x"0103060c",
  2048 => x"597f3e00",
  2049 => x"003e7f4d",
  2050 => x"7f060400",
  2051 => x"0000007f",
  2052 => x"71634200",
  2053 => x"00464f59",
  2054 => x"49632200",
  2055 => x"00367f49",
  2056 => x"13161c18",
  2057 => x"00107f7f",
  2058 => x"45672700",
  2059 => x"00397d45",
  2060 => x"4b7e3c00",
  2061 => x"00307949",
  2062 => x"71010100",
  2063 => x"00070f79",
  2064 => x"497f3600",
  2065 => x"00367f49",
  2066 => x"494f0600",
  2067 => x"001e3f69",
  2068 => x"66000000",
  2069 => x"00000066",
  2070 => x"e6800000",
  2071 => x"00000066",
  2072 => x"14080800",
  2073 => x"00222214",
  2074 => x"14141400",
  2075 => x"00141414",
  2076 => x"14222200",
  2077 => x"00080814",
  2078 => x"51030200",
  2079 => x"00060f59",
  2080 => x"5d417f3e",
  2081 => x"001e1f55",
  2082 => x"097f7e00",
  2083 => x"007e7f09",
  2084 => x"497f7f00",
  2085 => x"00367f49",
  2086 => x"633e1c00",
  2087 => x"00414141",
  2088 => x"417f7f00",
  2089 => x"001c3e63",
  2090 => x"497f7f00",
  2091 => x"00414149",
  2092 => x"097f7f00",
  2093 => x"00010109",
  2094 => x"417f3e00",
  2095 => x"007a7b49",
  2096 => x"087f7f00",
  2097 => x"007f7f08",
  2098 => x"7f410000",
  2099 => x"0000417f",
  2100 => x"40602000",
  2101 => x"003f7f40",
  2102 => x"1c087f7f",
  2103 => x"00416336",
  2104 => x"407f7f00",
  2105 => x"00404040",
  2106 => x"0c067f7f",
  2107 => x"007f7f06",
  2108 => x"0c067f7f",
  2109 => x"007f7f18",
  2110 => x"417f3e00",
  2111 => x"003e7f41",
  2112 => x"097f7f00",
  2113 => x"00060f09",
  2114 => x"61417f3e",
  2115 => x"00407e7f",
  2116 => x"097f7f00",
  2117 => x"00667f19",
  2118 => x"4d6f2600",
  2119 => x"00327b59",
  2120 => x"7f010100",
  2121 => x"0001017f",
  2122 => x"407f3f00",
  2123 => x"003f7f40",
  2124 => x"703f0f00",
  2125 => x"000f3f70",
  2126 => x"18307f7f",
  2127 => x"007f7f30",
  2128 => x"1c366341",
  2129 => x"4163361c",
  2130 => x"7c060301",
  2131 => x"0103067c",
  2132 => x"4d597161",
  2133 => x"00414347",
  2134 => x"7f7f0000",
  2135 => x"00004141",
  2136 => x"0c060301",
  2137 => x"40603018",
  2138 => x"41410000",
  2139 => x"00007f7f",
  2140 => x"03060c08",
  2141 => x"00080c06",
  2142 => x"80808080",
  2143 => x"00808080",
  2144 => x"03000000",
  2145 => x"00000407",
  2146 => x"54742000",
  2147 => x"00787c54",
  2148 => x"447f7f00",
  2149 => x"00387c44",
  2150 => x"447c3800",
  2151 => x"00004444",
  2152 => x"447c3800",
  2153 => x"007f7f44",
  2154 => x"547c3800",
  2155 => x"00185c54",
  2156 => x"7f7e0400",
  2157 => x"00000505",
  2158 => x"a4bc1800",
  2159 => x"007cfca4",
  2160 => x"047f7f00",
  2161 => x"00787c04",
  2162 => x"3d000000",
  2163 => x"0000407d",
  2164 => x"80808000",
  2165 => x"00007dfd",
  2166 => x"107f7f00",
  2167 => x"00446c38",
  2168 => x"3f000000",
  2169 => x"0000407f",
  2170 => x"180c7c7c",
  2171 => x"00787c0c",
  2172 => x"047c7c00",
  2173 => x"00787c04",
  2174 => x"447c3800",
  2175 => x"00387c44",
  2176 => x"24fcfc00",
  2177 => x"00183c24",
  2178 => x"243c1800",
  2179 => x"00fcfc24",
  2180 => x"047c7c00",
  2181 => x"00080c04",
  2182 => x"545c4800",
  2183 => x"00207454",
  2184 => x"7f3f0400",
  2185 => x"00004444",
  2186 => x"407c3c00",
  2187 => x"007c7c40",
  2188 => x"603c1c00",
  2189 => x"001c3c60",
  2190 => x"30607c3c",
  2191 => x"003c7c60",
  2192 => x"10386c44",
  2193 => x"00446c38",
  2194 => x"e0bc1c00",
  2195 => x"001c3c60",
  2196 => x"74644400",
  2197 => x"00444c5c",
  2198 => x"3e080800",
  2199 => x"00414177",
  2200 => x"7f000000",
  2201 => x"0000007f",
  2202 => x"77414100",
  2203 => x"0008083e",
  2204 => x"03010102",
  2205 => x"00010202",
  2206 => x"7f7f7f7f",
  2207 => x"007f7f7f",
  2208 => x"1c1c0808",
  2209 => x"7f7f3e3e",
  2210 => x"3e3e7f7f",
  2211 => x"08081c1c",
  2212 => x"7c181000",
  2213 => x"0010187c",
  2214 => x"7c301000",
  2215 => x"0010307c",
  2216 => x"60603010",
  2217 => x"00061e78",
  2218 => x"183c6642",
  2219 => x"0042663c",
  2220 => x"c26a3878",
  2221 => x"00386cc6",
  2222 => x"60000060",
  2223 => x"00600000",
  2224 => x"5c5b5e0e",
  2225 => x"86fc0e5d",
  2226 => x"f5c27e71",
  2227 => x"c04cbfd8",
  2228 => x"c41ec04b",
  2229 => x"c402ab66",
  2230 => x"c24dc087",
  2231 => x"754dc187",
  2232 => x"ee49731e",
  2233 => x"86c887e1",
  2234 => x"ef49e0c0",
  2235 => x"a4c487ea",
  2236 => x"f0496a4a",
  2237 => x"c8f187f1",
  2238 => x"c184cc87",
  2239 => x"abb7c883",
  2240 => x"87cdff04",
  2241 => x"4d268efc",
  2242 => x"4b264c26",
  2243 => x"711e4f26",
  2244 => x"dcf5c24a",
  2245 => x"dcf5c25a",
  2246 => x"4978c748",
  2247 => x"2687e1fe",
  2248 => x"1e731e4f",
  2249 => x"b7c04a71",
  2250 => x"87d303aa",
  2251 => x"bffcd9c2",
  2252 => x"c187c405",
  2253 => x"c087c24b",
  2254 => x"c0dac24b",
  2255 => x"c287c45b",
  2256 => x"fc5ac0da",
  2257 => x"fcd9c248",
  2258 => x"c14a78bf",
  2259 => x"a2c0c19a",
  2260 => x"87e6ec49",
  2261 => x"4f264b26",
  2262 => x"c44a711e",
  2263 => x"49721e66",
  2264 => x"fc87f0eb",
  2265 => x"1e4f268e",
  2266 => x"c348d4ff",
  2267 => x"d0ff78ff",
  2268 => x"78e1c048",
  2269 => x"c148d4ff",
  2270 => x"c4487178",
  2271 => x"08d4ff30",
  2272 => x"48d0ff78",
  2273 => x"2678e0c0",
  2274 => x"5b5e0e4f",
  2275 => x"ec0e5d5c",
  2276 => x"48a6c886",
  2277 => x"c47e78c0",
  2278 => x"78bfec80",
  2279 => x"f5c280f8",
  2280 => x"e878bfd8",
  2281 => x"d9c24cbf",
  2282 => x"e349bffc",
  2283 => x"eecb87eb",
  2284 => x"87cccb49",
  2285 => x"c758a6d4",
  2286 => x"87dfe749",
  2287 => x"c9059870",
  2288 => x"4966cc87",
  2289 => x"c10299c1",
  2290 => x"66d087c4",
  2291 => x"ec7ec14d",
  2292 => x"d9c24bbf",
  2293 => x"e249bffc",
  2294 => x"497587ff",
  2295 => x"7087edca",
  2296 => x"87d70298",
  2297 => x"bfe4d9c2",
  2298 => x"c2b9c149",
  2299 => x"7159e8d9",
  2300 => x"cb87f4fd",
  2301 => x"c7ca49ee",
  2302 => x"c74d7087",
  2303 => x"87dbe649",
  2304 => x"ff059870",
  2305 => x"497387c7",
  2306 => x"fe0599c1",
  2307 => x"026e87ff",
  2308 => x"c287e3c0",
  2309 => x"4abffcd9",
  2310 => x"dac2bac1",
  2311 => x"0afc5ac0",
  2312 => x"9ac10a7a",
  2313 => x"49a2c0c1",
  2314 => x"c187cfe9",
  2315 => x"eae549da",
  2316 => x"48a6c887",
  2317 => x"d9c278c1",
  2318 => x"c105bffc",
  2319 => x"c0c887c5",
  2320 => x"d9c24dc0",
  2321 => x"49134be8",
  2322 => x"87cfe549",
  2323 => x"c2029870",
  2324 => x"c1b47587",
  2325 => x"ff052db7",
  2326 => x"497487ec",
  2327 => x"7199ffc3",
  2328 => x"fb49c01e",
  2329 => x"497487f2",
  2330 => x"7129b7c8",
  2331 => x"fb49c11e",
  2332 => x"86c887e6",
  2333 => x"e449fdc3",
  2334 => x"fac387e1",
  2335 => x"87dbe449",
  2336 => x"7487d4c7",
  2337 => x"99ffc349",
  2338 => x"712cb7c8",
  2339 => x"029c74b4",
  2340 => x"d9c287df",
  2341 => x"c749bff8",
  2342 => x"987087f2",
  2343 => x"87c4c005",
  2344 => x"87d34cc0",
  2345 => x"c749e0c2",
  2346 => x"d9c287d6",
  2347 => x"c6c058fc",
  2348 => x"f8d9c287",
  2349 => x"7478c048",
  2350 => x"0599c849",
  2351 => x"c387cec0",
  2352 => x"d6e349f5",
  2353 => x"c2497087",
  2354 => x"e7c00299",
  2355 => x"dcf5c287",
  2356 => x"cac002bf",
  2357 => x"88c14887",
  2358 => x"58e0f5c2",
  2359 => x"c487d0c0",
  2360 => x"e0c14a66",
  2361 => x"c0026a82",
  2362 => x"ff4b87c5",
  2363 => x"c80f7349",
  2364 => x"78c148a6",
  2365 => x"99c44974",
  2366 => x"87cec005",
  2367 => x"e249f2c3",
  2368 => x"497087d9",
  2369 => x"c00299c2",
  2370 => x"f5c287f0",
  2371 => x"487ebfdc",
  2372 => x"03a8b7c7",
  2373 => x"6e87cbc0",
  2374 => x"c280c148",
  2375 => x"c058e0f5",
  2376 => x"66c487d3",
  2377 => x"80e0c148",
  2378 => x"bf6e7e70",
  2379 => x"87c5c002",
  2380 => x"7349fe4b",
  2381 => x"48a6c80f",
  2382 => x"fdc378c1",
  2383 => x"87dbe149",
  2384 => x"99c24970",
  2385 => x"87e9c002",
  2386 => x"bfdcf5c2",
  2387 => x"87c9c002",
  2388 => x"48dcf5c2",
  2389 => x"d3c078c0",
  2390 => x"4866c487",
  2391 => x"7080e0c1",
  2392 => x"02bf6e7e",
  2393 => x"4b87c5c0",
  2394 => x"0f7349fd",
  2395 => x"c148a6c8",
  2396 => x"49fac378",
  2397 => x"7087e4e0",
  2398 => x"0299c249",
  2399 => x"c287edc0",
  2400 => x"48bfdcf5",
  2401 => x"03a8b7c7",
  2402 => x"c287c9c0",
  2403 => x"c748dcf5",
  2404 => x"87d3c078",
  2405 => x"c14866c4",
  2406 => x"7e7080e0",
  2407 => x"c002bf6e",
  2408 => x"fc4b87c5",
  2409 => x"c80f7349",
  2410 => x"78c148a6",
  2411 => x"f5c27ec0",
  2412 => x"50c048d4",
  2413 => x"c349eecb",
  2414 => x"a6d487c6",
  2415 => x"d4f5c258",
  2416 => x"c105bf97",
  2417 => x"497487de",
  2418 => x"0599f0c3",
  2419 => x"c187cdc0",
  2420 => x"dfff49da",
  2421 => x"987087c5",
  2422 => x"87c8c102",
  2423 => x"bfe87ec1",
  2424 => x"ffc3494b",
  2425 => x"2bb7c899",
  2426 => x"d9c2b371",
  2427 => x"ff49bffc",
  2428 => x"d087e6da",
  2429 => x"d3c24966",
  2430 => x"02987087",
  2431 => x"c287c6c0",
  2432 => x"c148d4f5",
  2433 => x"d4f5c250",
  2434 => x"c005bf97",
  2435 => x"497387d6",
  2436 => x"0599f0c3",
  2437 => x"c187c5ff",
  2438 => x"ddff49da",
  2439 => x"987087fd",
  2440 => x"87f8fe05",
  2441 => x"e0c0026e",
  2442 => x"48a6cc87",
  2443 => x"bfdcf5c2",
  2444 => x"4966cc78",
  2445 => x"66c491cc",
  2446 => x"70807148",
  2447 => x"02bf6e7e",
  2448 => x"4b87c6c0",
  2449 => x"734966cc",
  2450 => x"0266c80f",
  2451 => x"c287c8c0",
  2452 => x"49bfdcf5",
  2453 => x"ec87e9f1",
  2454 => x"264d268e",
  2455 => x"264b264c",
  2456 => x"0000004f",
  2457 => x"00000000",
  2458 => x"14111258",
  2459 => x"231c1b1d",
  2460 => x"9491595a",
  2461 => x"f4ebf2f5",
  2462 => x"00000000",
  2463 => x"00000000",
  2464 => x"ff4a711e",
  2465 => x"7249bfc8",
  2466 => x"4f2648a1",
  2467 => x"bfc8ff1e",
  2468 => x"c0c0fe89",
  2469 => x"a9c0c0c0",
  2470 => x"c087c401",
  2471 => x"c187c24a",
  2472 => x"2648724a",
  2473 => x"5b5e0e4f",
  2474 => x"710e5d5c",
  2475 => x"4cd4ff4b",
  2476 => x"c04866d0",
  2477 => x"ff49d678",
  2478 => x"c387dddd",
  2479 => x"496c7cff",
  2480 => x"7199ffc3",
  2481 => x"f0c3494d",
  2482 => x"a9e0c199",
  2483 => x"c387cb05",
  2484 => x"486c7cff",
  2485 => x"66d098c3",
  2486 => x"ffc37808",
  2487 => x"494a6c7c",
  2488 => x"ffc331c8",
  2489 => x"714a6c7c",
  2490 => x"c84972b2",
  2491 => x"7cffc331",
  2492 => x"b2714a6c",
  2493 => x"31c84972",
  2494 => x"6c7cffc3",
  2495 => x"ffb2714a",
  2496 => x"e0c048d0",
  2497 => x"029b7378",
  2498 => x"7b7287c2",
  2499 => x"4d264875",
  2500 => x"4b264c26",
  2501 => x"261e4f26",
  2502 => x"5b5e0e4f",
  2503 => x"86f80e5c",
  2504 => x"a6c81e76",
  2505 => x"87fdfd49",
  2506 => x"4b7086c4",
  2507 => x"a8c2486e",
  2508 => x"87f0c203",
  2509 => x"f0c34a73",
  2510 => x"aad0c19a",
  2511 => x"c187c702",
  2512 => x"c205aae0",
  2513 => x"497387de",
  2514 => x"c30299c8",
  2515 => x"87c6ff87",
  2516 => x"9cc34c73",
  2517 => x"c105acc2",
  2518 => x"66c487c2",
  2519 => x"7131c949",
  2520 => x"4a66c41e",
  2521 => x"f5c292d4",
  2522 => x"817249e0",
  2523 => x"87e4cdfe",
  2524 => x"daff49d8",
  2525 => x"c0c887e2",
  2526 => x"f8e3c21e",
  2527 => x"d6e7fd49",
  2528 => x"48d0ff87",
  2529 => x"c278e0c0",
  2530 => x"cc1ef8e3",
  2531 => x"92d44a66",
  2532 => x"49e0f5c2",
  2533 => x"cbfe8172",
  2534 => x"86cc87eb",
  2535 => x"c105acc1",
  2536 => x"66c487c2",
  2537 => x"7131c949",
  2538 => x"4a66c41e",
  2539 => x"f5c292d4",
  2540 => x"817249e0",
  2541 => x"87dcccfe",
  2542 => x"1ef8e3c2",
  2543 => x"d44a66c8",
  2544 => x"e0f5c292",
  2545 => x"fe817249",
  2546 => x"d787ebc9",
  2547 => x"c7d9ff49",
  2548 => x"1ec0c887",
  2549 => x"49f8e3c2",
  2550 => x"87d8e5fd",
  2551 => x"d0ff86cc",
  2552 => x"78e0c048",
  2553 => x"4c268ef8",
  2554 => x"4f264b26",
  2555 => x"5c5b5e0e",
  2556 => x"86fc0e5d",
  2557 => x"d4ff4d71",
  2558 => x"7e66d44c",
  2559 => x"a8b7c348",
  2560 => x"87e2c101",
  2561 => x"66c41e75",
  2562 => x"c293d44b",
  2563 => x"7383e0f5",
  2564 => x"e0c3fe49",
  2565 => x"49a3c887",
  2566 => x"d0ff4969",
  2567 => x"78e1c848",
  2568 => x"48717cdd",
  2569 => x"7098ffc3",
  2570 => x"c84a717c",
  2571 => x"48722ab7",
  2572 => x"7098ffc3",
  2573 => x"d04a717c",
  2574 => x"48722ab7",
  2575 => x"7098ffc3",
  2576 => x"d848717c",
  2577 => x"7c7028b7",
  2578 => x"7c7c7cc0",
  2579 => x"7c7c7c7c",
  2580 => x"7c7c7c7c",
  2581 => x"48d0ff7c",
  2582 => x"c478e0c0",
  2583 => x"49dc1e66",
  2584 => x"87d9d7ff",
  2585 => x"8efc86c8",
  2586 => x"4c264d26",
  2587 => x"4f264b26",
  2588 => x"c01e731e",
  2589 => x"e2c21e4b",
  2590 => x"fd49bfec",
  2591 => x"86c487ee",
  2592 => x"bff0e2c2",
  2593 => x"fddbfe49",
  2594 => x"05987087",
  2595 => x"e2c287c4",
  2596 => x"48734bd8",
  2597 => x"4f264b26",
  2598 => x"204d4f52",
  2599 => x"64616f6c",
  2600 => x"20676e69",
  2601 => x"6c696166",
  2602 => x"00006465",
  2603 => x"000028b4",
  2604 => x"000028c0",
  2605 => x"20434242",
  2606 => x"20202020",
  2607 => x"00444856",
  2608 => x"20434242",
  2609 => x"20202020",
  2610 => x"004d4f52",
  2611 => x"00001baf",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
