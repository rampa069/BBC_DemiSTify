
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"59",x"7f",x"3e",x"00"),
     1 => (x"00",x"3e",x"7f",x"4d"),
     2 => (x"7f",x"06",x"04",x"00"),
     3 => (x"00",x"00",x"00",x"7f"),
     4 => (x"71",x"63",x"42",x"00"),
     5 => (x"00",x"46",x"4f",x"59"),
     6 => (x"49",x"63",x"22",x"00"),
     7 => (x"00",x"36",x"7f",x"49"),
     8 => (x"13",x"16",x"1c",x"18"),
     9 => (x"00",x"10",x"7f",x"7f"),
    10 => (x"45",x"67",x"27",x"00"),
    11 => (x"00",x"39",x"7d",x"45"),
    12 => (x"4b",x"7e",x"3c",x"00"),
    13 => (x"00",x"30",x"79",x"49"),
    14 => (x"71",x"01",x"01",x"00"),
    15 => (x"00",x"07",x"0f",x"79"),
    16 => (x"49",x"7f",x"36",x"00"),
    17 => (x"00",x"36",x"7f",x"49"),
    18 => (x"49",x"4f",x"06",x"00"),
    19 => (x"00",x"1e",x"3f",x"69"),
    20 => (x"66",x"00",x"00",x"00"),
    21 => (x"00",x"00",x"00",x"66"),
    22 => (x"e6",x"80",x"00",x"00"),
    23 => (x"00",x"00",x"00",x"66"),
    24 => (x"14",x"08",x"08",x"00"),
    25 => (x"00",x"22",x"22",x"14"),
    26 => (x"14",x"14",x"14",x"00"),
    27 => (x"00",x"14",x"14",x"14"),
    28 => (x"14",x"22",x"22",x"00"),
    29 => (x"00",x"08",x"08",x"14"),
    30 => (x"51",x"03",x"02",x"00"),
    31 => (x"00",x"06",x"0f",x"59"),
    32 => (x"5d",x"41",x"7f",x"3e"),
    33 => (x"00",x"1e",x"1f",x"55"),
    34 => (x"09",x"7f",x"7e",x"00"),
    35 => (x"00",x"7e",x"7f",x"09"),
    36 => (x"49",x"7f",x"7f",x"00"),
    37 => (x"00",x"36",x"7f",x"49"),
    38 => (x"63",x"3e",x"1c",x"00"),
    39 => (x"00",x"41",x"41",x"41"),
    40 => (x"41",x"7f",x"7f",x"00"),
    41 => (x"00",x"1c",x"3e",x"63"),
    42 => (x"49",x"7f",x"7f",x"00"),
    43 => (x"00",x"41",x"41",x"49"),
    44 => (x"09",x"7f",x"7f",x"00"),
    45 => (x"00",x"01",x"01",x"09"),
    46 => (x"41",x"7f",x"3e",x"00"),
    47 => (x"00",x"7a",x"7b",x"49"),
    48 => (x"08",x"7f",x"7f",x"00"),
    49 => (x"00",x"7f",x"7f",x"08"),
    50 => (x"7f",x"41",x"00",x"00"),
    51 => (x"00",x"00",x"41",x"7f"),
    52 => (x"40",x"60",x"20",x"00"),
    53 => (x"00",x"3f",x"7f",x"40"),
    54 => (x"1c",x"08",x"7f",x"7f"),
    55 => (x"00",x"41",x"63",x"36"),
    56 => (x"40",x"7f",x"7f",x"00"),
    57 => (x"00",x"40",x"40",x"40"),
    58 => (x"0c",x"06",x"7f",x"7f"),
    59 => (x"00",x"7f",x"7f",x"06"),
    60 => (x"0c",x"06",x"7f",x"7f"),
    61 => (x"00",x"7f",x"7f",x"18"),
    62 => (x"41",x"7f",x"3e",x"00"),
    63 => (x"00",x"3e",x"7f",x"41"),
    64 => (x"09",x"7f",x"7f",x"00"),
    65 => (x"00",x"06",x"0f",x"09"),
    66 => (x"61",x"41",x"7f",x"3e"),
    67 => (x"00",x"40",x"7e",x"7f"),
    68 => (x"09",x"7f",x"7f",x"00"),
    69 => (x"00",x"66",x"7f",x"19"),
    70 => (x"4d",x"6f",x"26",x"00"),
    71 => (x"00",x"32",x"7b",x"59"),
    72 => (x"7f",x"01",x"01",x"00"),
    73 => (x"00",x"01",x"01",x"7f"),
    74 => (x"40",x"7f",x"3f",x"00"),
    75 => (x"00",x"3f",x"7f",x"40"),
    76 => (x"70",x"3f",x"0f",x"00"),
    77 => (x"00",x"0f",x"3f",x"70"),
    78 => (x"18",x"30",x"7f",x"7f"),
    79 => (x"00",x"7f",x"7f",x"30"),
    80 => (x"1c",x"36",x"63",x"41"),
    81 => (x"41",x"63",x"36",x"1c"),
    82 => (x"7c",x"06",x"03",x"01"),
    83 => (x"01",x"03",x"06",x"7c"),
    84 => (x"4d",x"59",x"71",x"61"),
    85 => (x"00",x"41",x"43",x"47"),
    86 => (x"7f",x"7f",x"00",x"00"),
    87 => (x"00",x"00",x"41",x"41"),
    88 => (x"0c",x"06",x"03",x"01"),
    89 => (x"40",x"60",x"30",x"18"),
    90 => (x"41",x"41",x"00",x"00"),
    91 => (x"00",x"00",x"7f",x"7f"),
    92 => (x"03",x"06",x"0c",x"08"),
    93 => (x"00",x"08",x"0c",x"06"),
    94 => (x"80",x"80",x"80",x"80"),
    95 => (x"00",x"80",x"80",x"80"),
    96 => (x"03",x"00",x"00",x"00"),
    97 => (x"00",x"00",x"04",x"07"),
    98 => (x"54",x"74",x"20",x"00"),
    99 => (x"00",x"78",x"7c",x"54"),
   100 => (x"44",x"7f",x"7f",x"00"),
   101 => (x"00",x"38",x"7c",x"44"),
   102 => (x"44",x"7c",x"38",x"00"),
   103 => (x"00",x"00",x"44",x"44"),
   104 => (x"44",x"7c",x"38",x"00"),
   105 => (x"00",x"7f",x"7f",x"44"),
   106 => (x"54",x"7c",x"38",x"00"),
   107 => (x"00",x"18",x"5c",x"54"),
   108 => (x"7f",x"7e",x"04",x"00"),
   109 => (x"00",x"00",x"05",x"05"),
   110 => (x"a4",x"bc",x"18",x"00"),
   111 => (x"00",x"7c",x"fc",x"a4"),
   112 => (x"04",x"7f",x"7f",x"00"),
   113 => (x"00",x"78",x"7c",x"04"),
   114 => (x"3d",x"00",x"00",x"00"),
   115 => (x"00",x"00",x"40",x"7d"),
   116 => (x"80",x"80",x"80",x"00"),
   117 => (x"00",x"00",x"7d",x"fd"),
   118 => (x"10",x"7f",x"7f",x"00"),
   119 => (x"00",x"44",x"6c",x"38"),
   120 => (x"3f",x"00",x"00",x"00"),
   121 => (x"00",x"00",x"40",x"7f"),
   122 => (x"18",x"0c",x"7c",x"7c"),
   123 => (x"00",x"78",x"7c",x"0c"),
   124 => (x"04",x"7c",x"7c",x"00"),
   125 => (x"00",x"78",x"7c",x"04"),
   126 => (x"44",x"7c",x"38",x"00"),
   127 => (x"00",x"38",x"7c",x"44"),
   128 => (x"24",x"fc",x"fc",x"00"),
   129 => (x"00",x"18",x"3c",x"24"),
   130 => (x"24",x"3c",x"18",x"00"),
   131 => (x"00",x"fc",x"fc",x"24"),
   132 => (x"04",x"7c",x"7c",x"00"),
   133 => (x"00",x"08",x"0c",x"04"),
   134 => (x"54",x"5c",x"48",x"00"),
   135 => (x"00",x"20",x"74",x"54"),
   136 => (x"7f",x"3f",x"04",x"00"),
   137 => (x"00",x"00",x"44",x"44"),
   138 => (x"40",x"7c",x"3c",x"00"),
   139 => (x"00",x"7c",x"7c",x"40"),
   140 => (x"60",x"3c",x"1c",x"00"),
   141 => (x"00",x"1c",x"3c",x"60"),
   142 => (x"30",x"60",x"7c",x"3c"),
   143 => (x"00",x"3c",x"7c",x"60"),
   144 => (x"10",x"38",x"6c",x"44"),
   145 => (x"00",x"44",x"6c",x"38"),
   146 => (x"e0",x"bc",x"1c",x"00"),
   147 => (x"00",x"1c",x"3c",x"60"),
   148 => (x"74",x"64",x"44",x"00"),
   149 => (x"00",x"44",x"4c",x"5c"),
   150 => (x"3e",x"08",x"08",x"00"),
   151 => (x"00",x"41",x"41",x"77"),
   152 => (x"7f",x"00",x"00",x"00"),
   153 => (x"00",x"00",x"00",x"7f"),
   154 => (x"77",x"41",x"41",x"00"),
   155 => (x"00",x"08",x"08",x"3e"),
   156 => (x"03",x"01",x"01",x"02"),
   157 => (x"00",x"01",x"02",x"02"),
   158 => (x"7f",x"7f",x"7f",x"7f"),
   159 => (x"00",x"7f",x"7f",x"7f"),
   160 => (x"1c",x"1c",x"08",x"08"),
   161 => (x"7f",x"7f",x"3e",x"3e"),
   162 => (x"3e",x"3e",x"7f",x"7f"),
   163 => (x"08",x"08",x"1c",x"1c"),
   164 => (x"7c",x"18",x"10",x"00"),
   165 => (x"00",x"10",x"18",x"7c"),
   166 => (x"7c",x"30",x"10",x"00"),
   167 => (x"00",x"10",x"30",x"7c"),
   168 => (x"60",x"60",x"30",x"10"),
   169 => (x"00",x"06",x"1e",x"78"),
   170 => (x"18",x"3c",x"66",x"42"),
   171 => (x"00",x"42",x"66",x"3c"),
   172 => (x"c2",x"6a",x"38",x"78"),
   173 => (x"00",x"38",x"6c",x"c6"),
   174 => (x"60",x"00",x"00",x"60"),
   175 => (x"00",x"60",x"00",x"00"),
   176 => (x"5c",x"5b",x"5e",x"0e"),
   177 => (x"86",x"fc",x"0e",x"5d"),
   178 => (x"f5",x"c2",x"7e",x"71"),
   179 => (x"c0",x"4c",x"bf",x"d8"),
   180 => (x"c4",x"1e",x"c0",x"4b"),
   181 => (x"c4",x"02",x"ab",x"66"),
   182 => (x"c2",x"4d",x"c0",x"87"),
   183 => (x"75",x"4d",x"c1",x"87"),
   184 => (x"ee",x"49",x"73",x"1e"),
   185 => (x"86",x"c8",x"87",x"e1"),
   186 => (x"ef",x"49",x"e0",x"c0"),
   187 => (x"a4",x"c4",x"87",x"ea"),
   188 => (x"f0",x"49",x"6a",x"4a"),
   189 => (x"c8",x"f1",x"87",x"f1"),
   190 => (x"c1",x"84",x"cc",x"87"),
   191 => (x"ab",x"b7",x"c8",x"83"),
   192 => (x"87",x"cd",x"ff",x"04"),
   193 => (x"4d",x"26",x"8e",x"fc"),
   194 => (x"4b",x"26",x"4c",x"26"),
   195 => (x"71",x"1e",x"4f",x"26"),
   196 => (x"dc",x"f5",x"c2",x"4a"),
   197 => (x"dc",x"f5",x"c2",x"5a"),
   198 => (x"49",x"78",x"c7",x"48"),
   199 => (x"26",x"87",x"e1",x"fe"),
   200 => (x"1e",x"73",x"1e",x"4f"),
   201 => (x"b7",x"c0",x"4a",x"71"),
   202 => (x"87",x"d3",x"03",x"aa"),
   203 => (x"bf",x"fc",x"d9",x"c2"),
   204 => (x"c1",x"87",x"c4",x"05"),
   205 => (x"c0",x"87",x"c2",x"4b"),
   206 => (x"c0",x"da",x"c2",x"4b"),
   207 => (x"c2",x"87",x"c4",x"5b"),
   208 => (x"fc",x"5a",x"c0",x"da"),
   209 => (x"fc",x"d9",x"c2",x"48"),
   210 => (x"c1",x"4a",x"78",x"bf"),
   211 => (x"a2",x"c0",x"c1",x"9a"),
   212 => (x"87",x"e6",x"ec",x"49"),
   213 => (x"4f",x"26",x"4b",x"26"),
   214 => (x"c4",x"4a",x"71",x"1e"),
   215 => (x"49",x"72",x"1e",x"66"),
   216 => (x"fc",x"87",x"f0",x"eb"),
   217 => (x"1e",x"4f",x"26",x"8e"),
   218 => (x"c3",x"48",x"d4",x"ff"),
   219 => (x"d0",x"ff",x"78",x"ff"),
   220 => (x"78",x"e1",x"c0",x"48"),
   221 => (x"c1",x"48",x"d4",x"ff"),
   222 => (x"c4",x"48",x"71",x"78"),
   223 => (x"08",x"d4",x"ff",x"30"),
   224 => (x"48",x"d0",x"ff",x"78"),
   225 => (x"26",x"78",x"e0",x"c0"),
   226 => (x"5b",x"5e",x"0e",x"4f"),
   227 => (x"ec",x"0e",x"5d",x"5c"),
   228 => (x"48",x"a6",x"c8",x"86"),
   229 => (x"c4",x"7e",x"78",x"c0"),
   230 => (x"78",x"bf",x"ec",x"80"),
   231 => (x"f5",x"c2",x"80",x"f8"),
   232 => (x"e8",x"78",x"bf",x"d8"),
   233 => (x"d9",x"c2",x"4c",x"bf"),
   234 => (x"e3",x"49",x"bf",x"fc"),
   235 => (x"ee",x"cb",x"87",x"eb"),
   236 => (x"87",x"cc",x"cb",x"49"),
   237 => (x"c7",x"58",x"a6",x"d4"),
   238 => (x"87",x"df",x"e7",x"49"),
   239 => (x"c9",x"05",x"98",x"70"),
   240 => (x"49",x"66",x"cc",x"87"),
   241 => (x"c1",x"02",x"99",x"c1"),
   242 => (x"66",x"d0",x"87",x"c4"),
   243 => (x"ec",x"7e",x"c1",x"4d"),
   244 => (x"d9",x"c2",x"4b",x"bf"),
   245 => (x"e2",x"49",x"bf",x"fc"),
   246 => (x"49",x"75",x"87",x"ff"),
   247 => (x"70",x"87",x"ed",x"ca"),
   248 => (x"87",x"d7",x"02",x"98"),
   249 => (x"bf",x"e4",x"d9",x"c2"),
   250 => (x"c2",x"b9",x"c1",x"49"),
   251 => (x"71",x"59",x"e8",x"d9"),
   252 => (x"cb",x"87",x"f4",x"fd"),
   253 => (x"c7",x"ca",x"49",x"ee"),
   254 => (x"c7",x"4d",x"70",x"87"),
   255 => (x"87",x"db",x"e6",x"49"),
   256 => (x"ff",x"05",x"98",x"70"),
   257 => (x"49",x"73",x"87",x"c7"),
   258 => (x"fe",x"05",x"99",x"c1"),
   259 => (x"02",x"6e",x"87",x"ff"),
   260 => (x"c2",x"87",x"e3",x"c0"),
   261 => (x"4a",x"bf",x"fc",x"d9"),
   262 => (x"da",x"c2",x"ba",x"c1"),
   263 => (x"0a",x"fc",x"5a",x"c0"),
   264 => (x"9a",x"c1",x"0a",x"7a"),
   265 => (x"49",x"a2",x"c0",x"c1"),
   266 => (x"c1",x"87",x"cf",x"e9"),
   267 => (x"ea",x"e5",x"49",x"da"),
   268 => (x"48",x"a6",x"c8",x"87"),
   269 => (x"d9",x"c2",x"78",x"c1"),
   270 => (x"c1",x"05",x"bf",x"fc"),
   271 => (x"c0",x"c8",x"87",x"c5"),
   272 => (x"d9",x"c2",x"4d",x"c0"),
   273 => (x"49",x"13",x"4b",x"e8"),
   274 => (x"87",x"cf",x"e5",x"49"),
   275 => (x"c2",x"02",x"98",x"70"),
   276 => (x"c1",x"b4",x"75",x"87"),
   277 => (x"ff",x"05",x"2d",x"b7"),
   278 => (x"49",x"74",x"87",x"ec"),
   279 => (x"71",x"99",x"ff",x"c3"),
   280 => (x"fb",x"49",x"c0",x"1e"),
   281 => (x"49",x"74",x"87",x"f2"),
   282 => (x"71",x"29",x"b7",x"c8"),
   283 => (x"fb",x"49",x"c1",x"1e"),
   284 => (x"86",x"c8",x"87",x"e6"),
   285 => (x"e4",x"49",x"fd",x"c3"),
   286 => (x"fa",x"c3",x"87",x"e1"),
   287 => (x"87",x"db",x"e4",x"49"),
   288 => (x"74",x"87",x"d4",x"c7"),
   289 => (x"99",x"ff",x"c3",x"49"),
   290 => (x"71",x"2c",x"b7",x"c8"),
   291 => (x"02",x"9c",x"74",x"b4"),
   292 => (x"d9",x"c2",x"87",x"df"),
   293 => (x"c7",x"49",x"bf",x"f8"),
   294 => (x"98",x"70",x"87",x"f2"),
   295 => (x"87",x"c4",x"c0",x"05"),
   296 => (x"87",x"d3",x"4c",x"c0"),
   297 => (x"c7",x"49",x"e0",x"c2"),
   298 => (x"d9",x"c2",x"87",x"d6"),
   299 => (x"c6",x"c0",x"58",x"fc"),
   300 => (x"f8",x"d9",x"c2",x"87"),
   301 => (x"74",x"78",x"c0",x"48"),
   302 => (x"05",x"99",x"c8",x"49"),
   303 => (x"c3",x"87",x"ce",x"c0"),
   304 => (x"d6",x"e3",x"49",x"f5"),
   305 => (x"c2",x"49",x"70",x"87"),
   306 => (x"e7",x"c0",x"02",x"99"),
   307 => (x"dc",x"f5",x"c2",x"87"),
   308 => (x"ca",x"c0",x"02",x"bf"),
   309 => (x"88",x"c1",x"48",x"87"),
   310 => (x"58",x"e0",x"f5",x"c2"),
   311 => (x"c4",x"87",x"d0",x"c0"),
   312 => (x"e0",x"c1",x"4a",x"66"),
   313 => (x"c0",x"02",x"6a",x"82"),
   314 => (x"ff",x"4b",x"87",x"c5"),
   315 => (x"c8",x"0f",x"73",x"49"),
   316 => (x"78",x"c1",x"48",x"a6"),
   317 => (x"99",x"c4",x"49",x"74"),
   318 => (x"87",x"ce",x"c0",x"05"),
   319 => (x"e2",x"49",x"f2",x"c3"),
   320 => (x"49",x"70",x"87",x"d9"),
   321 => (x"c0",x"02",x"99",x"c2"),
   322 => (x"f5",x"c2",x"87",x"f0"),
   323 => (x"48",x"7e",x"bf",x"dc"),
   324 => (x"03",x"a8",x"b7",x"c7"),
   325 => (x"6e",x"87",x"cb",x"c0"),
   326 => (x"c2",x"80",x"c1",x"48"),
   327 => (x"c0",x"58",x"e0",x"f5"),
   328 => (x"66",x"c4",x"87",x"d3"),
   329 => (x"80",x"e0",x"c1",x"48"),
   330 => (x"bf",x"6e",x"7e",x"70"),
   331 => (x"87",x"c5",x"c0",x"02"),
   332 => (x"73",x"49",x"fe",x"4b"),
   333 => (x"48",x"a6",x"c8",x"0f"),
   334 => (x"fd",x"c3",x"78",x"c1"),
   335 => (x"87",x"db",x"e1",x"49"),
   336 => (x"99",x"c2",x"49",x"70"),
   337 => (x"87",x"e9",x"c0",x"02"),
   338 => (x"bf",x"dc",x"f5",x"c2"),
   339 => (x"87",x"c9",x"c0",x"02"),
   340 => (x"48",x"dc",x"f5",x"c2"),
   341 => (x"d3",x"c0",x"78",x"c0"),
   342 => (x"48",x"66",x"c4",x"87"),
   343 => (x"70",x"80",x"e0",x"c1"),
   344 => (x"02",x"bf",x"6e",x"7e"),
   345 => (x"4b",x"87",x"c5",x"c0"),
   346 => (x"0f",x"73",x"49",x"fd"),
   347 => (x"c1",x"48",x"a6",x"c8"),
   348 => (x"49",x"fa",x"c3",x"78"),
   349 => (x"70",x"87",x"e4",x"e0"),
   350 => (x"02",x"99",x"c2",x"49"),
   351 => (x"c2",x"87",x"ed",x"c0"),
   352 => (x"48",x"bf",x"dc",x"f5"),
   353 => (x"03",x"a8",x"b7",x"c7"),
   354 => (x"c2",x"87",x"c9",x"c0"),
   355 => (x"c7",x"48",x"dc",x"f5"),
   356 => (x"87",x"d3",x"c0",x"78"),
   357 => (x"c1",x"48",x"66",x"c4"),
   358 => (x"7e",x"70",x"80",x"e0"),
   359 => (x"c0",x"02",x"bf",x"6e"),
   360 => (x"fc",x"4b",x"87",x"c5"),
   361 => (x"c8",x"0f",x"73",x"49"),
   362 => (x"78",x"c1",x"48",x"a6"),
   363 => (x"f5",x"c2",x"7e",x"c0"),
   364 => (x"50",x"c0",x"48",x"d4"),
   365 => (x"c3",x"49",x"ee",x"cb"),
   366 => (x"a6",x"d4",x"87",x"c6"),
   367 => (x"d4",x"f5",x"c2",x"58"),
   368 => (x"c1",x"05",x"bf",x"97"),
   369 => (x"49",x"74",x"87",x"de"),
   370 => (x"05",x"99",x"f0",x"c3"),
   371 => (x"c1",x"87",x"cd",x"c0"),
   372 => (x"df",x"ff",x"49",x"da"),
   373 => (x"98",x"70",x"87",x"c5"),
   374 => (x"87",x"c8",x"c1",x"02"),
   375 => (x"bf",x"e8",x"7e",x"c1"),
   376 => (x"ff",x"c3",x"49",x"4b"),
   377 => (x"2b",x"b7",x"c8",x"99"),
   378 => (x"d9",x"c2",x"b3",x"71"),
   379 => (x"ff",x"49",x"bf",x"fc"),
   380 => (x"d0",x"87",x"e6",x"da"),
   381 => (x"d3",x"c2",x"49",x"66"),
   382 => (x"02",x"98",x"70",x"87"),
   383 => (x"c2",x"87",x"c6",x"c0"),
   384 => (x"c1",x"48",x"d4",x"f5"),
   385 => (x"d4",x"f5",x"c2",x"50"),
   386 => (x"c0",x"05",x"bf",x"97"),
   387 => (x"49",x"73",x"87",x"d6"),
   388 => (x"05",x"99",x"f0",x"c3"),
   389 => (x"c1",x"87",x"c5",x"ff"),
   390 => (x"dd",x"ff",x"49",x"da"),
   391 => (x"98",x"70",x"87",x"fd"),
   392 => (x"87",x"f8",x"fe",x"05"),
   393 => (x"e0",x"c0",x"02",x"6e"),
   394 => (x"48",x"a6",x"cc",x"87"),
   395 => (x"bf",x"dc",x"f5",x"c2"),
   396 => (x"49",x"66",x"cc",x"78"),
   397 => (x"66",x"c4",x"91",x"cc"),
   398 => (x"70",x"80",x"71",x"48"),
   399 => (x"02",x"bf",x"6e",x"7e"),
   400 => (x"4b",x"87",x"c6",x"c0"),
   401 => (x"73",x"49",x"66",x"cc"),
   402 => (x"02",x"66",x"c8",x"0f"),
   403 => (x"c2",x"87",x"c8",x"c0"),
   404 => (x"49",x"bf",x"dc",x"f5"),
   405 => (x"ec",x"87",x"e9",x"f1"),
   406 => (x"26",x"4d",x"26",x"8e"),
   407 => (x"26",x"4b",x"26",x"4c"),
   408 => (x"00",x"00",x"00",x"4f"),
   409 => (x"00",x"00",x"00",x"00"),
   410 => (x"14",x"11",x"12",x"58"),
   411 => (x"23",x"1c",x"1b",x"1d"),
   412 => (x"94",x"91",x"59",x"5a"),
   413 => (x"f4",x"eb",x"f2",x"f5"),
   414 => (x"00",x"00",x"00",x"00"),
   415 => (x"00",x"00",x"00",x"00"),
   416 => (x"ff",x"4a",x"71",x"1e"),
   417 => (x"72",x"49",x"bf",x"c8"),
   418 => (x"4f",x"26",x"48",x"a1"),
   419 => (x"bf",x"c8",x"ff",x"1e"),
   420 => (x"c0",x"c0",x"fe",x"89"),
   421 => (x"a9",x"c0",x"c0",x"c0"),
   422 => (x"c0",x"87",x"c4",x"01"),
   423 => (x"c1",x"87",x"c2",x"4a"),
   424 => (x"26",x"48",x"72",x"4a"),
   425 => (x"5b",x"5e",x"0e",x"4f"),
   426 => (x"71",x"0e",x"5d",x"5c"),
   427 => (x"4c",x"d4",x"ff",x"4b"),
   428 => (x"c0",x"48",x"66",x"d0"),
   429 => (x"ff",x"49",x"d6",x"78"),
   430 => (x"c3",x"87",x"dd",x"dd"),
   431 => (x"49",x"6c",x"7c",x"ff"),
   432 => (x"71",x"99",x"ff",x"c3"),
   433 => (x"f0",x"c3",x"49",x"4d"),
   434 => (x"a9",x"e0",x"c1",x"99"),
   435 => (x"c3",x"87",x"cb",x"05"),
   436 => (x"48",x"6c",x"7c",x"ff"),
   437 => (x"66",x"d0",x"98",x"c3"),
   438 => (x"ff",x"c3",x"78",x"08"),
   439 => (x"49",x"4a",x"6c",x"7c"),
   440 => (x"ff",x"c3",x"31",x"c8"),
   441 => (x"71",x"4a",x"6c",x"7c"),
   442 => (x"c8",x"49",x"72",x"b2"),
   443 => (x"7c",x"ff",x"c3",x"31"),
   444 => (x"b2",x"71",x"4a",x"6c"),
   445 => (x"31",x"c8",x"49",x"72"),
   446 => (x"6c",x"7c",x"ff",x"c3"),
   447 => (x"ff",x"b2",x"71",x"4a"),
   448 => (x"e0",x"c0",x"48",x"d0"),
   449 => (x"02",x"9b",x"73",x"78"),
   450 => (x"7b",x"72",x"87",x"c2"),
   451 => (x"4d",x"26",x"48",x"75"),
   452 => (x"4b",x"26",x"4c",x"26"),
   453 => (x"26",x"1e",x"4f",x"26"),
   454 => (x"5b",x"5e",x"0e",x"4f"),
   455 => (x"86",x"f8",x"0e",x"5c"),
   456 => (x"a6",x"c8",x"1e",x"76"),
   457 => (x"87",x"fd",x"fd",x"49"),
   458 => (x"4b",x"70",x"86",x"c4"),
   459 => (x"a8",x"c2",x"48",x"6e"),
   460 => (x"87",x"f0",x"c2",x"03"),
   461 => (x"f0",x"c3",x"4a",x"73"),
   462 => (x"aa",x"d0",x"c1",x"9a"),
   463 => (x"c1",x"87",x"c7",x"02"),
   464 => (x"c2",x"05",x"aa",x"e0"),
   465 => (x"49",x"73",x"87",x"de"),
   466 => (x"c3",x"02",x"99",x"c8"),
   467 => (x"87",x"c6",x"ff",x"87"),
   468 => (x"9c",x"c3",x"4c",x"73"),
   469 => (x"c1",x"05",x"ac",x"c2"),
   470 => (x"66",x"c4",x"87",x"c2"),
   471 => (x"71",x"31",x"c9",x"49"),
   472 => (x"4a",x"66",x"c4",x"1e"),
   473 => (x"f5",x"c2",x"92",x"d4"),
   474 => (x"81",x"72",x"49",x"e0"),
   475 => (x"87",x"e4",x"cd",x"fe"),
   476 => (x"da",x"ff",x"49",x"d8"),
   477 => (x"c0",x"c8",x"87",x"e2"),
   478 => (x"f8",x"e3",x"c2",x"1e"),
   479 => (x"d6",x"e7",x"fd",x"49"),
   480 => (x"48",x"d0",x"ff",x"87"),
   481 => (x"c2",x"78",x"e0",x"c0"),
   482 => (x"cc",x"1e",x"f8",x"e3"),
   483 => (x"92",x"d4",x"4a",x"66"),
   484 => (x"49",x"e0",x"f5",x"c2"),
   485 => (x"cb",x"fe",x"81",x"72"),
   486 => (x"86",x"cc",x"87",x"eb"),
   487 => (x"c1",x"05",x"ac",x"c1"),
   488 => (x"66",x"c4",x"87",x"c2"),
   489 => (x"71",x"31",x"c9",x"49"),
   490 => (x"4a",x"66",x"c4",x"1e"),
   491 => (x"f5",x"c2",x"92",x"d4"),
   492 => (x"81",x"72",x"49",x"e0"),
   493 => (x"87",x"dc",x"cc",x"fe"),
   494 => (x"1e",x"f8",x"e3",x"c2"),
   495 => (x"d4",x"4a",x"66",x"c8"),
   496 => (x"e0",x"f5",x"c2",x"92"),
   497 => (x"fe",x"81",x"72",x"49"),
   498 => (x"d7",x"87",x"eb",x"c9"),
   499 => (x"c7",x"d9",x"ff",x"49"),
   500 => (x"1e",x"c0",x"c8",x"87"),
   501 => (x"49",x"f8",x"e3",x"c2"),
   502 => (x"87",x"d8",x"e5",x"fd"),
   503 => (x"d0",x"ff",x"86",x"cc"),
   504 => (x"78",x"e0",x"c0",x"48"),
   505 => (x"4c",x"26",x"8e",x"f8"),
   506 => (x"4f",x"26",x"4b",x"26"),
   507 => (x"5c",x"5b",x"5e",x"0e"),
   508 => (x"86",x"fc",x"0e",x"5d"),
   509 => (x"d4",x"ff",x"4d",x"71"),
   510 => (x"7e",x"66",x"d4",x"4c"),
   511 => (x"a8",x"b7",x"c3",x"48"),
   512 => (x"87",x"e2",x"c1",x"01"),
   513 => (x"66",x"c4",x"1e",x"75"),
   514 => (x"c2",x"93",x"d4",x"4b"),
   515 => (x"73",x"83",x"e0",x"f5"),
   516 => (x"e0",x"c3",x"fe",x"49"),
   517 => (x"49",x"a3",x"c8",x"87"),
   518 => (x"d0",x"ff",x"49",x"69"),
   519 => (x"78",x"e1",x"c8",x"48"),
   520 => (x"48",x"71",x"7c",x"dd"),
   521 => (x"70",x"98",x"ff",x"c3"),
   522 => (x"c8",x"4a",x"71",x"7c"),
   523 => (x"48",x"72",x"2a",x"b7"),
   524 => (x"70",x"98",x"ff",x"c3"),
   525 => (x"d0",x"4a",x"71",x"7c"),
   526 => (x"48",x"72",x"2a",x"b7"),
   527 => (x"70",x"98",x"ff",x"c3"),
   528 => (x"d8",x"48",x"71",x"7c"),
   529 => (x"7c",x"70",x"28",x"b7"),
   530 => (x"7c",x"7c",x"7c",x"c0"),
   531 => (x"7c",x"7c",x"7c",x"7c"),
   532 => (x"7c",x"7c",x"7c",x"7c"),
   533 => (x"48",x"d0",x"ff",x"7c"),
   534 => (x"c4",x"78",x"e0",x"c0"),
   535 => (x"49",x"dc",x"1e",x"66"),
   536 => (x"87",x"d9",x"d7",x"ff"),
   537 => (x"8e",x"fc",x"86",x"c8"),
   538 => (x"4c",x"26",x"4d",x"26"),
   539 => (x"4f",x"26",x"4b",x"26"),
   540 => (x"c0",x"1e",x"73",x"1e"),
   541 => (x"e2",x"c2",x"1e",x"4b"),
   542 => (x"fd",x"49",x"bf",x"ec"),
   543 => (x"86",x"c4",x"87",x"ee"),
   544 => (x"bf",x"f0",x"e2",x"c2"),
   545 => (x"fd",x"db",x"fe",x"49"),
   546 => (x"05",x"98",x"70",x"87"),
   547 => (x"e2",x"c2",x"87",x"c4"),
   548 => (x"48",x"73",x"4b",x"d8"),
   549 => (x"4f",x"26",x"4b",x"26"),
   550 => (x"20",x"4d",x"4f",x"52"),
   551 => (x"64",x"61",x"6f",x"6c"),
   552 => (x"20",x"67",x"6e",x"69"),
   553 => (x"6c",x"69",x"61",x"66"),
   554 => (x"00",x"00",x"64",x"65"),
   555 => (x"00",x"00",x"28",x"b4"),
   556 => (x"00",x"00",x"28",x"c0"),
   557 => (x"20",x"43",x"42",x"42"),
   558 => (x"20",x"20",x"20",x"20"),
   559 => (x"00",x"44",x"48",x"56"),
   560 => (x"20",x"43",x"42",x"42"),
   561 => (x"20",x"20",x"20",x"20"),
   562 => (x"00",x"4d",x"4f",x"52"),
   563 => (x"00",x"00",x"1b",x"af"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

