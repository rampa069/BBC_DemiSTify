library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c4f6c287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49c4f6c2",
    18 => x"48cce3c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"cce3c287",
    25 => x"c8e3c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e8c187f7",
    29 => x"e3c287c2",
    30 => x"e3c24dcc",
    31 => x"ad744ccc",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"731e741e",
    65 => x"c11e721e",
    66 => x"87d0048b",
    67 => x"02114812",
    68 => x"c34c87ca",
    69 => x"749c98df",
    70 => x"87eb0288",
    71 => x"4b264a26",
    72 => x"4f264c26",
    73 => x"8148731e",
    74 => x"c502a973",
    75 => x"05531287",
    76 => x"4f2687f6",
    77 => x"711e731e",
    78 => x"4b66c84a",
    79 => x"718bc149",
    80 => x"87cf0299",
    81 => x"d4ff4812",
    82 => x"49737808",
    83 => x"99718bc1",
    84 => x"2687f105",
    85 => x"0e4f264b",
    86 => x"0e5c5b5e",
    87 => x"d4ff4a71",
    88 => x"4b66cc4c",
    89 => x"718bc149",
    90 => x"87ce0299",
    91 => x"6c7cffc3",
    92 => x"c1497352",
    93 => x"0599718b",
    94 => x"4c2687f2",
    95 => x"4f264b26",
    96 => x"ff1e731e",
    97 => x"ffc34bd4",
    98 => x"c34a6b7b",
    99 => x"496b7bff",
   100 => x"b17232c8",
   101 => x"6b7bffc3",
   102 => x"7131c84a",
   103 => x"7bffc3b2",
   104 => x"32c8496b",
   105 => x"4871b172",
   106 => x"4f264b26",
   107 => x"5c5b5e0e",
   108 => x"4d710e5d",
   109 => x"754cd4ff",
   110 => x"98ffc348",
   111 => x"e3c27c70",
   112 => x"c805bfcc",
   113 => x"4866d087",
   114 => x"a6d430c9",
   115 => x"4966d058",
   116 => x"487129d8",
   117 => x"7098ffc3",
   118 => x"4966d07c",
   119 => x"487129d0",
   120 => x"7098ffc3",
   121 => x"4966d07c",
   122 => x"487129c8",
   123 => x"7098ffc3",
   124 => x"4866d07c",
   125 => x"7098ffc3",
   126 => x"d049757c",
   127 => x"c3487129",
   128 => x"7c7098ff",
   129 => x"f0c94b6c",
   130 => x"ffc34aff",
   131 => x"87cf05ab",
   132 => x"6c7c7149",
   133 => x"028ac14b",
   134 => x"ab7187c5",
   135 => x"7387f202",
   136 => x"264d2648",
   137 => x"264b264c",
   138 => x"49c01e4f",
   139 => x"c348d4ff",
   140 => x"81c178ff",
   141 => x"a9b7c8c3",
   142 => x"2687f104",
   143 => x"5b5e0e4f",
   144 => x"c00e5d5c",
   145 => x"f7c1f0ff",
   146 => x"c0c0c14d",
   147 => x"4bc0c0c0",
   148 => x"c487d6ff",
   149 => x"c04cdff8",
   150 => x"fd49751e",
   151 => x"86c487ce",
   152 => x"c005a8c1",
   153 => x"d4ff87e5",
   154 => x"78ffc348",
   155 => x"e1c01e73",
   156 => x"49e9c1f0",
   157 => x"c487f5fc",
   158 => x"05987086",
   159 => x"d4ff87ca",
   160 => x"78ffc348",
   161 => x"87cb48c1",
   162 => x"c187defe",
   163 => x"c6ff058c",
   164 => x"2648c087",
   165 => x"264c264d",
   166 => x"0e4f264b",
   167 => x"0e5c5b5e",
   168 => x"c1f0ffc0",
   169 => x"d4ff4cc1",
   170 => x"78ffc348",
   171 => x"f749e0cb",
   172 => x"4bd387f5",
   173 => x"49741ec0",
   174 => x"c487f1fb",
   175 => x"05987086",
   176 => x"d4ff87ca",
   177 => x"78ffc348",
   178 => x"87cb48c1",
   179 => x"c187dafd",
   180 => x"dfff058b",
   181 => x"2648c087",
   182 => x"264b264c",
   183 => x"0000004f",
   184 => x"00444d43",
   185 => x"5c5b5e0e",
   186 => x"ffc30e5d",
   187 => x"4bd4ff4d",
   188 => x"c687f6fc",
   189 => x"e1c01eea",
   190 => x"49c8c1f0",
   191 => x"c487edfa",
   192 => x"02a8c186",
   193 => x"d2fe87c8",
   194 => x"c148c087",
   195 => x"eff987e8",
   196 => x"cf497087",
   197 => x"c699ffff",
   198 => x"c802a9ea",
   199 => x"87fbfd87",
   200 => x"d1c148c0",
   201 => x"c07b7587",
   202 => x"d0fc4cf1",
   203 => x"02987087",
   204 => x"c087ecc0",
   205 => x"f0ffc01e",
   206 => x"f949fac1",
   207 => x"86c487ee",
   208 => x"da059870",
   209 => x"6b7b7587",
   210 => x"757b7549",
   211 => x"757b757b",
   212 => x"99c0c17b",
   213 => x"c187c402",
   214 => x"c087db48",
   215 => x"c287d748",
   216 => x"87ca05ac",
   217 => x"f449c0ce",
   218 => x"48c087fd",
   219 => x"8cc187c8",
   220 => x"87f6fe05",
   221 => x"4d2648c0",
   222 => x"4b264c26",
   223 => x"00004f26",
   224 => x"43484453",
   225 => x"69616620",
   226 => x"000a216c",
   227 => x"5c5b5e0e",
   228 => x"d0ff0e5d",
   229 => x"d0e5c04d",
   230 => x"c24cc0c1",
   231 => x"c148cce3",
   232 => x"49d8d078",
   233 => x"c787c0f4",
   234 => x"f97dc24b",
   235 => x"7dc387fb",
   236 => x"49741ec0",
   237 => x"c487f5f7",
   238 => x"05a8c186",
   239 => x"c24b87c1",
   240 => x"87cb05ab",
   241 => x"f349d0d0",
   242 => x"48c087dd",
   243 => x"c187f6c0",
   244 => x"d4ff058b",
   245 => x"87ccfc87",
   246 => x"58d0e3c2",
   247 => x"cd059870",
   248 => x"c01ec187",
   249 => x"d0c1f0ff",
   250 => x"87c0f749",
   251 => x"d4ff86c4",
   252 => x"78ffc348",
   253 => x"c287ccc5",
   254 => x"c258d4e3",
   255 => x"48d4ff7d",
   256 => x"c178ffc3",
   257 => x"264d2648",
   258 => x"264b264c",
   259 => x"0000004f",
   260 => x"52524549",
   261 => x"00000000",
   262 => x"00495053",
   263 => x"5c5b5e0e",
   264 => x"4d710e5d",
   265 => x"ff4cffc3",
   266 => x"7b744bd4",
   267 => x"c448d0ff",
   268 => x"7b7478c3",
   269 => x"ffc01e75",
   270 => x"49d8c1f0",
   271 => x"c487edf5",
   272 => x"02987086",
   273 => x"c8d287cb",
   274 => x"87dbf149",
   275 => x"eec048c1",
   276 => x"c37b7487",
   277 => x"c0c87bfe",
   278 => x"4966d41e",
   279 => x"c487d5f3",
   280 => x"747b7486",
   281 => x"d87b747b",
   282 => x"744ae0da",
   283 => x"c5056b7b",
   284 => x"058ac187",
   285 => x"7b7487f5",
   286 => x"c248d0ff",
   287 => x"2648c078",
   288 => x"264c264d",
   289 => x"004f264b",
   290 => x"74697257",
   291 => x"61662065",
   292 => x"64656c69",
   293 => x"5e0e000a",
   294 => x"0e5d5c5b",
   295 => x"4b7186fc",
   296 => x"c04cd4ff",
   297 => x"cdeec57e",
   298 => x"ffc34adf",
   299 => x"c3486c7c",
   300 => x"c005a8fe",
   301 => x"4d7487f8",
   302 => x"cc029b73",
   303 => x"1e66d487",
   304 => x"d2f24973",
   305 => x"d486c487",
   306 => x"48d0ff87",
   307 => x"d478d1c4",
   308 => x"ffc34a66",
   309 => x"058ac17d",
   310 => x"a6d887f8",
   311 => x"7cffc35a",
   312 => x"059b737c",
   313 => x"d0ff87c5",
   314 => x"c178d048",
   315 => x"8ac17e4a",
   316 => x"87f6fe05",
   317 => x"8efc486e",
   318 => x"4c264d26",
   319 => x"4f264b26",
   320 => x"711e731e",
   321 => x"ff4bc04a",
   322 => x"ffc348d4",
   323 => x"48d0ff78",
   324 => x"ff78c3c4",
   325 => x"ffc348d4",
   326 => x"c01e7278",
   327 => x"d1c1f0ff",
   328 => x"87c8f249",
   329 => x"987086c4",
   330 => x"c887d205",
   331 => x"66cc1ec0",
   332 => x"87e2fd49",
   333 => x"4b7086c4",
   334 => x"c248d0ff",
   335 => x"26487378",
   336 => x"0e4f264b",
   337 => x"5d5c5b5e",
   338 => x"c01ec00e",
   339 => x"c9c1f0ff",
   340 => x"87d8f149",
   341 => x"e3c21ed2",
   342 => x"f9fc49d4",
   343 => x"c086c887",
   344 => x"d284c14c",
   345 => x"f804acb7",
   346 => x"d4e3c287",
   347 => x"c349bf97",
   348 => x"c0c199c0",
   349 => x"e7c005a9",
   350 => x"dbe3c287",
   351 => x"d049bf97",
   352 => x"dce3c231",
   353 => x"c84abf97",
   354 => x"c2b17232",
   355 => x"bf97dde3",
   356 => x"4c71b14a",
   357 => x"ffffffcf",
   358 => x"ca84c19c",
   359 => x"87e7c134",
   360 => x"97dde3c2",
   361 => x"31c149bf",
   362 => x"e3c299c6",
   363 => x"4abf97de",
   364 => x"722ab7c7",
   365 => x"d9e3c2b1",
   366 => x"4d4abf97",
   367 => x"e3c29dcf",
   368 => x"4abf97da",
   369 => x"32ca9ac3",
   370 => x"97dbe3c2",
   371 => x"33c24bbf",
   372 => x"e3c2b273",
   373 => x"4bbf97dc",
   374 => x"c69bc0c3",
   375 => x"b2732bb7",
   376 => x"48c181c2",
   377 => x"49703071",
   378 => x"307548c1",
   379 => x"4c724d70",
   380 => x"947184c1",
   381 => x"adb7c0c8",
   382 => x"c187cc06",
   383 => x"c82db734",
   384 => x"01adb7c0",
   385 => x"7487f4ff",
   386 => x"264d2648",
   387 => x"264b264c",
   388 => x"5b5e0e4f",
   389 => x"f80e5d5c",
   390 => x"fcebc286",
   391 => x"c278c048",
   392 => x"c01ef4e3",
   393 => x"87d8fb49",
   394 => x"987086c4",
   395 => x"c087c505",
   396 => x"87c0c948",
   397 => x"7ec14dc0",
   398 => x"bfd8f7c0",
   399 => x"eae4c249",
   400 => x"4bc8714a",
   401 => x"7087dfea",
   402 => x"87c20598",
   403 => x"f7c07ec0",
   404 => x"c249bfd4",
   405 => x"714ac6e5",
   406 => x"c9ea4bc8",
   407 => x"05987087",
   408 => x"7ec087c2",
   409 => x"fdc0026e",
   410 => x"faeac287",
   411 => x"ebc24dbf",
   412 => x"7ebf9ff2",
   413 => x"ead6c548",
   414 => x"87c705a8",
   415 => x"bffaeac2",
   416 => x"6e87ce4d",
   417 => x"d5e9ca48",
   418 => x"87c502a8",
   419 => x"e3c748c0",
   420 => x"f4e3c287",
   421 => x"f949751e",
   422 => x"86c487e6",
   423 => x"c5059870",
   424 => x"c748c087",
   425 => x"f7c087ce",
   426 => x"c249bfd4",
   427 => x"714ac6e5",
   428 => x"f1e84bc8",
   429 => x"05987087",
   430 => x"ebc287c8",
   431 => x"78c148fc",
   432 => x"f7c087da",
   433 => x"c249bfd8",
   434 => x"714aeae4",
   435 => x"d5e84bc8",
   436 => x"02987087",
   437 => x"c087c5c0",
   438 => x"87d8c648",
   439 => x"97f2ebc2",
   440 => x"d5c149bf",
   441 => x"cdc005a9",
   442 => x"f3ebc287",
   443 => x"c249bf97",
   444 => x"c002a9ea",
   445 => x"48c087c5",
   446 => x"c287f9c5",
   447 => x"bf97f4e3",
   448 => x"e9c3487e",
   449 => x"cec002a8",
   450 => x"c3486e87",
   451 => x"c002a8eb",
   452 => x"48c087c5",
   453 => x"c287ddc5",
   454 => x"bf97ffe3",
   455 => x"c0059949",
   456 => x"e4c287cc",
   457 => x"49bf97c0",
   458 => x"c002a9c2",
   459 => x"48c087c5",
   460 => x"c287c1c5",
   461 => x"bf97c1e4",
   462 => x"f8ebc248",
   463 => x"484c7058",
   464 => x"ebc288c1",
   465 => x"e4c258fc",
   466 => x"49bf97c2",
   467 => x"e4c28175",
   468 => x"4abf97c3",
   469 => x"a17232c8",
   470 => x"ccf0c27e",
   471 => x"c2786e48",
   472 => x"bf97c4e4",
   473 => x"58a6c848",
   474 => x"bffcebc2",
   475 => x"87cfc202",
   476 => x"bfd4f7c0",
   477 => x"c6e5c249",
   478 => x"4bc8714a",
   479 => x"7087e7e5",
   480 => x"c5c00298",
   481 => x"c348c087",
   482 => x"ebc287ea",
   483 => x"c24cbff4",
   484 => x"c25ce0f0",
   485 => x"bf97d9e4",
   486 => x"c231c849",
   487 => x"bf97d8e4",
   488 => x"c249a14a",
   489 => x"bf97dae4",
   490 => x"7232d04a",
   491 => x"e4c249a1",
   492 => x"4abf97db",
   493 => x"a17232d8",
   494 => x"9166c449",
   495 => x"bfccf0c2",
   496 => x"d4f0c281",
   497 => x"e1e4c259",
   498 => x"c84abf97",
   499 => x"e0e4c232",
   500 => x"a24bbf97",
   501 => x"e2e4c24a",
   502 => x"d04bbf97",
   503 => x"4aa27333",
   504 => x"97e3e4c2",
   505 => x"9bcf4bbf",
   506 => x"a27333d8",
   507 => x"d8f0c24a",
   508 => x"748ac25a",
   509 => x"d8f0c292",
   510 => x"78a17248",
   511 => x"c287c1c1",
   512 => x"bf97c6e4",
   513 => x"c231c849",
   514 => x"bf97c5e4",
   515 => x"c549a14a",
   516 => x"81ffc731",
   517 => x"f0c229c9",
   518 => x"e4c259e0",
   519 => x"4abf97cb",
   520 => x"e4c232c8",
   521 => x"4bbf97ca",
   522 => x"66c44aa2",
   523 => x"c2826e92",
   524 => x"c25adcf0",
   525 => x"c048d4f0",
   526 => x"d0f0c278",
   527 => x"78a17248",
   528 => x"48e0f0c2",
   529 => x"bfd4f0c2",
   530 => x"e4f0c278",
   531 => x"d8f0c248",
   532 => x"ebc278bf",
   533 => x"c002bffc",
   534 => x"487487c9",
   535 => x"7e7030c4",
   536 => x"c287c9c0",
   537 => x"48bfdcf0",
   538 => x"7e7030c4",
   539 => x"48c0ecc2",
   540 => x"48c1786e",
   541 => x"4d268ef8",
   542 => x"4b264c26",
   543 => x"5e0e4f26",
   544 => x"0e5d5c5b",
   545 => x"ebc24a71",
   546 => x"cb02bffc",
   547 => x"c74b7287",
   548 => x"c14d722b",
   549 => x"87c99dff",
   550 => x"2bc84b72",
   551 => x"ffc34d72",
   552 => x"ccf0c29d",
   553 => x"f7c083bf",
   554 => x"02abbfd0",
   555 => x"f7c087d9",
   556 => x"e3c25bd4",
   557 => x"49731ef4",
   558 => x"c487c5f1",
   559 => x"05987086",
   560 => x"48c087c5",
   561 => x"c287e6c0",
   562 => x"02bffceb",
   563 => x"497587d2",
   564 => x"e3c291c4",
   565 => x"4c6981f4",
   566 => x"ffffffcf",
   567 => x"87cb9cff",
   568 => x"91c24975",
   569 => x"81f4e3c2",
   570 => x"744c699f",
   571 => x"264d2648",
   572 => x"264b264c",
   573 => x"5b5e0e4f",
   574 => x"f40e5d5c",
   575 => x"59a6cc86",
   576 => x"c50566c8",
   577 => x"c348c087",
   578 => x"66c887c7",
   579 => x"7080c848",
   580 => x"78c0487e",
   581 => x"c70266dc",
   582 => x"9766dc87",
   583 => x"87c505bf",
   584 => x"ecc248c0",
   585 => x"c11ec087",
   586 => x"e9ca4949",
   587 => x"7086c487",
   588 => x"c0029c4c",
   589 => x"ecc287fc",
   590 => x"66dc4ac4",
   591 => x"cadeff49",
   592 => x"02987087",
   593 => x"7487ebc0",
   594 => x"4966dc4a",
   595 => x"deff4bcb",
   596 => x"987087ee",
   597 => x"c087db02",
   598 => x"029c741e",
   599 => x"4dc087c4",
   600 => x"4dc187c2",
   601 => x"edc94975",
   602 => x"7086c487",
   603 => x"ff059c4c",
   604 => x"9c7487c4",
   605 => x"87d7c102",
   606 => x"6e49a4dc",
   607 => x"da786948",
   608 => x"66c849a4",
   609 => x"c880c448",
   610 => x"699f58a6",
   611 => x"0866c448",
   612 => x"fcebc278",
   613 => x"87d202bf",
   614 => x"9f49a4d4",
   615 => x"ffc04969",
   616 => x"487199ff",
   617 => x"7e7030d0",
   618 => x"7ec087c2",
   619 => x"66c4486e",
   620 => x"66c480bf",
   621 => x"66c87808",
   622 => x"c878c048",
   623 => x"81cc4966",
   624 => x"79bf66c4",
   625 => x"d04966c8",
   626 => x"c179c081",
   627 => x"c087c248",
   628 => x"268ef448",
   629 => x"264c264d",
   630 => x"0e4f264b",
   631 => x"5d5c5b5e",
   632 => x"d04c710e",
   633 => x"9c744d66",
   634 => x"87c2c102",
   635 => x"6949a4c8",
   636 => x"87fac002",
   637 => x"7585496c",
   638 => x"f8ebc2b9",
   639 => x"baff4abf",
   640 => x"99719972",
   641 => x"87e4c002",
   642 => x"6b4ba4c4",
   643 => x"87eef949",
   644 => x"ebc27b70",
   645 => x"6c49bff4",
   646 => x"757c7181",
   647 => x"f8ebc2b9",
   648 => x"baff4abf",
   649 => x"99719972",
   650 => x"87dcff05",
   651 => x"4d267c75",
   652 => x"4b264c26",
   653 => x"731e4f26",
   654 => x"9b4b711e",
   655 => x"c887c702",
   656 => x"056949a3",
   657 => x"48c087c5",
   658 => x"c287f6c0",
   659 => x"49bfd0f0",
   660 => x"6a4aa3c4",
   661 => x"c28ac24a",
   662 => x"92bff4eb",
   663 => x"c249a172",
   664 => x"4abff8eb",
   665 => x"a1729a6b",
   666 => x"d4f7c049",
   667 => x"1e66c859",
   668 => x"87ccea71",
   669 => x"987086c4",
   670 => x"c087c405",
   671 => x"c187c248",
   672 => x"264b2648",
   673 => x"1e731e4f",
   674 => x"029b4b71",
   675 => x"a3c887c7",
   676 => x"c5056949",
   677 => x"c048c087",
   678 => x"f0c287f6",
   679 => x"c449bfd0",
   680 => x"4a6a4aa3",
   681 => x"ebc28ac2",
   682 => x"7292bff4",
   683 => x"ebc249a1",
   684 => x"6b4abff8",
   685 => x"49a1729a",
   686 => x"59d4f7c0",
   687 => x"711e66c8",
   688 => x"c487d9e5",
   689 => x"05987086",
   690 => x"48c087c4",
   691 => x"48c187c2",
   692 => x"4f264b26",
   693 => x"5c5b5e0e",
   694 => x"86fc0e5d",
   695 => x"66d44b71",
   696 => x"029b734d",
   697 => x"c887ccc1",
   698 => x"026949a3",
   699 => x"d087c4c1",
   700 => x"ebc24ca3",
   701 => x"ff49bff8",
   702 => x"994a6cb9",
   703 => x"a966d47e",
   704 => x"c087cd06",
   705 => x"a3cc7c7b",
   706 => x"49a3c44a",
   707 => x"87ca796a",
   708 => x"c0f84972",
   709 => x"4d66d499",
   710 => x"49758d71",
   711 => x"1e7129c9",
   712 => x"f6fa4973",
   713 => x"f4e3c287",
   714 => x"fc49731e",
   715 => x"86c887c8",
   716 => x"fc7c66d4",
   717 => x"264d268e",
   718 => x"264b264c",
   719 => x"1e731e4f",
   720 => x"029b4b71",
   721 => x"c287e4c0",
   722 => x"735be4f0",
   723 => x"c28ac24a",
   724 => x"49bff4eb",
   725 => x"d0f0c292",
   726 => x"807248bf",
   727 => x"58e8f0c2",
   728 => x"30c44871",
   729 => x"58c4ecc2",
   730 => x"c287edc0",
   731 => x"c248e0f0",
   732 => x"78bfd4f0",
   733 => x"48e4f0c2",
   734 => x"bfd8f0c2",
   735 => x"fcebc278",
   736 => x"87c902bf",
   737 => x"bff4ebc2",
   738 => x"c731c449",
   739 => x"dcf0c287",
   740 => x"31c449bf",
   741 => x"59c4ecc2",
   742 => x"4f264b26",
   743 => x"5c5b5e0e",
   744 => x"c04a710e",
   745 => x"029a724b",
   746 => x"da87e0c0",
   747 => x"699f49a2",
   748 => x"fcebc24b",
   749 => x"87cf02bf",
   750 => x"9f49a2d4",
   751 => x"c04c4969",
   752 => x"d09cffff",
   753 => x"c087c234",
   754 => x"73b3744c",
   755 => x"87edfd49",
   756 => x"4b264c26",
   757 => x"5e0e4f26",
   758 => x"0e5d5c5b",
   759 => x"a6c886f0",
   760 => x"ffffcf59",
   761 => x"c04cf8ff",
   762 => x"0266c47e",
   763 => x"e3c287d8",
   764 => x"78c048f0",
   765 => x"48e8e3c2",
   766 => x"bfe4f0c2",
   767 => x"ece3c278",
   768 => x"e0f0c248",
   769 => x"ecc278bf",
   770 => x"50c048d1",
   771 => x"bfc0ecc2",
   772 => x"f0e3c249",
   773 => x"aa714abf",
   774 => x"87cbc403",
   775 => x"99cf4972",
   776 => x"87e9c005",
   777 => x"48d0f7c0",
   778 => x"bfe8e3c2",
   779 => x"f4e3c278",
   780 => x"e8e3c21e",
   781 => x"e3c249bf",
   782 => x"a1c148e8",
   783 => x"ffe27178",
   784 => x"c086c487",
   785 => x"c248ccf7",
   786 => x"cc78f4e3",
   787 => x"ccf7c087",
   788 => x"e0c048bf",
   789 => x"d0f7c080",
   790 => x"f0e3c258",
   791 => x"80c148bf",
   792 => x"58f4e3c2",
   793 => x"000dcc27",
   794 => x"bf97bf00",
   795 => x"c2029d4d",
   796 => x"e5c387e5",
   797 => x"dec202ad",
   798 => x"ccf7c087",
   799 => x"a3cb4bbf",
   800 => x"cf4c1149",
   801 => x"d2c105ac",
   802 => x"df497587",
   803 => x"cd89c199",
   804 => x"c4ecc291",
   805 => x"4aa3c181",
   806 => x"a3c35112",
   807 => x"c551124a",
   808 => x"51124aa3",
   809 => x"124aa3c7",
   810 => x"4aa3c951",
   811 => x"a3ce5112",
   812 => x"d051124a",
   813 => x"51124aa3",
   814 => x"124aa3d2",
   815 => x"4aa3d451",
   816 => x"a3d65112",
   817 => x"d851124a",
   818 => x"51124aa3",
   819 => x"124aa3dc",
   820 => x"4aa3de51",
   821 => x"7ec15112",
   822 => x"7487fcc0",
   823 => x"0599c849",
   824 => x"7487edc0",
   825 => x"0599d049",
   826 => x"e0c087d3",
   827 => x"ccc00266",
   828 => x"c0497387",
   829 => x"700f66e0",
   830 => x"d3c00298",
   831 => x"c0056e87",
   832 => x"ecc287c6",
   833 => x"50c048c4",
   834 => x"bfccf7c0",
   835 => x"87e9c248",
   836 => x"48d1ecc2",
   837 => x"c27e50c0",
   838 => x"49bfc0ec",
   839 => x"bff0e3c2",
   840 => x"04aa714a",
   841 => x"cf87f5fb",
   842 => x"f8ffffff",
   843 => x"e4f0c24c",
   844 => x"c8c005bf",
   845 => x"fcebc287",
   846 => x"fac102bf",
   847 => x"ece3c287",
   848 => x"f9ec49bf",
   849 => x"f0e3c287",
   850 => x"48a6c458",
   851 => x"bfece3c2",
   852 => x"fcebc278",
   853 => x"dbc002bf",
   854 => x"4966c487",
   855 => x"a9749974",
   856 => x"87c8c002",
   857 => x"c048a6c8",
   858 => x"87e7c078",
   859 => x"c148a6c8",
   860 => x"87dfc078",
   861 => x"cf4966c4",
   862 => x"a999f8ff",
   863 => x"87c8c002",
   864 => x"c048a6cc",
   865 => x"87c5c078",
   866 => x"c148a6cc",
   867 => x"48a6c878",
   868 => x"c87866cc",
   869 => x"dec00566",
   870 => x"4966c487",
   871 => x"ebc289c2",
   872 => x"c291bff4",
   873 => x"48bfd0f0",
   874 => x"e3c28071",
   875 => x"e3c258ec",
   876 => x"78c048f0",
   877 => x"c087d5f9",
   878 => x"ffffcf48",
   879 => x"f04cf8ff",
   880 => x"264d268e",
   881 => x"264b264c",
   882 => x"0000004f",
   883 => x"00000000",
   884 => x"ffffffff",
   885 => x"00000ddc",
   886 => x"00000de8",
   887 => x"33544146",
   888 => x"20202032",
   889 => x"00000000",
   890 => x"31544146",
   891 => x"20202036",
   892 => x"d4ff1e00",
   893 => x"78ffc348",
   894 => x"4f264868",
   895 => x"48d4ff1e",
   896 => x"ff78ffc3",
   897 => x"e1c048d0",
   898 => x"48d4ff78",
   899 => x"4f2678d4",
   900 => x"48d0ff1e",
   901 => x"2678e0c0",
   902 => x"d4ff1e4f",
   903 => x"99497087",
   904 => x"c087c602",
   905 => x"f105a9fb",
   906 => x"26487187",
   907 => x"5b5e0e4f",
   908 => x"4b710e5c",
   909 => x"f8fe4cc0",
   910 => x"99497087",
   911 => x"87f9c002",
   912 => x"02a9ecc0",
   913 => x"c087f2c0",
   914 => x"c002a9fb",
   915 => x"66cc87eb",
   916 => x"c703acb7",
   917 => x"0266d087",
   918 => x"537187c2",
   919 => x"c2029971",
   920 => x"fe84c187",
   921 => x"497087cb",
   922 => x"87cd0299",
   923 => x"02a9ecc0",
   924 => x"fbc087c7",
   925 => x"d5ff05a9",
   926 => x"0266d087",
   927 => x"97c087c3",
   928 => x"a9ecc07b",
   929 => x"7487c405",
   930 => x"7487c54a",
   931 => x"8a0ac04a",
   932 => x"4c264872",
   933 => x"4f264b26",
   934 => x"87d5fd1e",
   935 => x"c04a4970",
   936 => x"c904aaf0",
   937 => x"aaf9c087",
   938 => x"c087c301",
   939 => x"c1c18af0",
   940 => x"87c904aa",
   941 => x"01aadac1",
   942 => x"f7c087c3",
   943 => x"2648728a",
   944 => x"5b5e0e4f",
   945 => x"f80e5d5c",
   946 => x"c04c7186",
   947 => x"87ecfc7e",
   948 => x"fdc04bc0",
   949 => x"49bf97e0",
   950 => x"cf04a9c0",
   951 => x"87f9fc87",
   952 => x"fdc083c1",
   953 => x"49bf97e0",
   954 => x"87f106ab",
   955 => x"97e0fdc0",
   956 => x"87cf02bf",
   957 => x"7087fafb",
   958 => x"c6029949",
   959 => x"a9ecc087",
   960 => x"c087f105",
   961 => x"87e9fb4b",
   962 => x"e4fb4d70",
   963 => x"58a6c887",
   964 => x"7087defb",
   965 => x"c883c14a",
   966 => x"699749a4",
   967 => x"da05ad49",
   968 => x"49a4c987",
   969 => x"c4496997",
   970 => x"ce05a966",
   971 => x"49a4ca87",
   972 => x"aa496997",
   973 => x"c187c405",
   974 => x"c087d07e",
   975 => x"c602adec",
   976 => x"adfbc087",
   977 => x"c087c405",
   978 => x"6e7ec14b",
   979 => x"87f5fe02",
   980 => x"7387fdfa",
   981 => x"268ef848",
   982 => x"264c264d",
   983 => x"004f264b",
   984 => x"1e731e00",
   985 => x"c84bd4ff",
   986 => x"d0ff4a66",
   987 => x"78c5c848",
   988 => x"c148d4ff",
   989 => x"7b1178d4",
   990 => x"f9058ac1",
   991 => x"48d0ff87",
   992 => x"4b2678c4",
   993 => x"5e0e4f26",
   994 => x"0e5d5c5b",
   995 => x"7e7186f8",
   996 => x"f0c21e6e",
   997 => x"dce549f4",
   998 => x"7086c487",
   999 => x"e4c40298",
  1000 => x"e4ecc187",
  1001 => x"496e4cbf",
  1002 => x"c887d6fc",
  1003 => x"987058a6",
  1004 => x"c487c505",
  1005 => x"78c148a6",
  1006 => x"c548d0ff",
  1007 => x"48d4ff78",
  1008 => x"c478d5c1",
  1009 => x"89c14966",
  1010 => x"ecc131c6",
  1011 => x"4abf97dc",
  1012 => x"ffb07148",
  1013 => x"ff7808d4",
  1014 => x"78c448d0",
  1015 => x"97f0f0c2",
  1016 => x"99d049bf",
  1017 => x"c587dd02",
  1018 => x"48d4ff78",
  1019 => x"c078d6c1",
  1020 => x"48d4ff4a",
  1021 => x"c178ffc3",
  1022 => x"aae0c082",
  1023 => x"ff87f204",
  1024 => x"78c448d0",
  1025 => x"c348d4ff",
  1026 => x"d0ff78ff",
  1027 => x"ff78c548",
  1028 => x"d3c148d4",
  1029 => x"ff78c178",
  1030 => x"78c448d0",
  1031 => x"06acb7c0",
  1032 => x"c287cbc2",
  1033 => x"4bbffcf0",
  1034 => x"737e748c",
  1035 => x"ddc1029b",
  1036 => x"4dc0c887",
  1037 => x"abb7c08b",
  1038 => x"c887c603",
  1039 => x"c04da3c0",
  1040 => x"f0f0c24b",
  1041 => x"d049bf97",
  1042 => x"87cf0299",
  1043 => x"f0c21ec0",
  1044 => x"e1e749f4",
  1045 => x"7086c487",
  1046 => x"c287d84c",
  1047 => x"c21ef4e3",
  1048 => x"e749f4f0",
  1049 => x"4c7087d0",
  1050 => x"e3c21e75",
  1051 => x"f0fb49f4",
  1052 => x"7486c887",
  1053 => x"87c5059c",
  1054 => x"cac148c0",
  1055 => x"c21ec187",
  1056 => x"e549f4f0",
  1057 => x"86c487d5",
  1058 => x"fe059b73",
  1059 => x"4c6e87e3",
  1060 => x"06acb7c0",
  1061 => x"f0c287d1",
  1062 => x"78c048f4",
  1063 => x"78c080d0",
  1064 => x"f1c280f4",
  1065 => x"c078bfc0",
  1066 => x"fd01acb7",
  1067 => x"d0ff87f5",
  1068 => x"ff78c548",
  1069 => x"d3c148d4",
  1070 => x"ff78c078",
  1071 => x"78c448d0",
  1072 => x"c2c048c1",
  1073 => x"f848c087",
  1074 => x"264d268e",
  1075 => x"264b264c",
  1076 => x"5b5e0e4f",
  1077 => x"fc0e5d5c",
  1078 => x"c04d7186",
  1079 => x"04ad4c4b",
  1080 => x"c087e8c0",
  1081 => x"741ec1fb",
  1082 => x"87c4029c",
  1083 => x"87c24ac0",
  1084 => x"49724ac1",
  1085 => x"c487dfeb",
  1086 => x"c17e7086",
  1087 => x"c2056e83",
  1088 => x"c14b7587",
  1089 => x"06ab7584",
  1090 => x"6e87d8ff",
  1091 => x"268efc48",
  1092 => x"264c264d",
  1093 => x"0e4f264b",
  1094 => x"0e5c5b5e",
  1095 => x"66cc4b71",
  1096 => x"4c87d802",
  1097 => x"028cf0c0",
  1098 => x"4a7487d8",
  1099 => x"d1028ac1",
  1100 => x"cd028a87",
  1101 => x"c9028a87",
  1102 => x"7387d987",
  1103 => x"87c6f949",
  1104 => x"1e7487d2",
  1105 => x"dac149c0",
  1106 => x"1e7487de",
  1107 => x"dac14973",
  1108 => x"86c887d6",
  1109 => x"4b264c26",
  1110 => x"5e0e4f26",
  1111 => x"0e5d5c5b",
  1112 => x"4c7186fc",
  1113 => x"c291de49",
  1114 => x"714de0f1",
  1115 => x"026d9785",
  1116 => x"c287dcc1",
  1117 => x"49bfd0f1",
  1118 => x"fd718174",
  1119 => x"7e7087d3",
  1120 => x"c0029848",
  1121 => x"f1c287f2",
  1122 => x"4a704bd4",
  1123 => x"fefe49cb",
  1124 => x"4b7487d2",
  1125 => x"ecc193cc",
  1126 => x"83c483e8",
  1127 => x"7bdcc7c1",
  1128 => x"c4c14974",
  1129 => x"7b7587d6",
  1130 => x"97e0ecc1",
  1131 => x"c21e49bf",
  1132 => x"fd49d4f1",
  1133 => x"86c487e1",
  1134 => x"c3c14974",
  1135 => x"49c087fe",
  1136 => x"87d9c5c1",
  1137 => x"48ecf0c2",
  1138 => x"c04950c0",
  1139 => x"fc87c8e2",
  1140 => x"264d268e",
  1141 => x"264b264c",
  1142 => x"0000004f",
  1143 => x"64616f4c",
  1144 => x"2e676e69",
  1145 => x"1e002e2e",
  1146 => x"4b711e73",
  1147 => x"d0f1c249",
  1148 => x"fb7181bf",
  1149 => x"4a7087db",
  1150 => x"87c4029a",
  1151 => x"87dce649",
  1152 => x"48d0f1c2",
  1153 => x"497378c0",
  1154 => x"2687fac1",
  1155 => x"1e4f264b",
  1156 => x"4b711e73",
  1157 => x"024aa3c4",
  1158 => x"c187d0c1",
  1159 => x"87dc028a",
  1160 => x"f2c0028a",
  1161 => x"c1058a87",
  1162 => x"f1c287d3",
  1163 => x"c102bfd0",
  1164 => x"c14887cb",
  1165 => x"d4f1c288",
  1166 => x"87c1c158",
  1167 => x"bfd0f1c2",
  1168 => x"c289c649",
  1169 => x"c059d4f1",
  1170 => x"c003a9b7",
  1171 => x"f1c287ef",
  1172 => x"78c048d0",
  1173 => x"c287e6c0",
  1174 => x"02bfccf1",
  1175 => x"f1c287df",
  1176 => x"c148bfd0",
  1177 => x"d4f1c280",
  1178 => x"c287d258",
  1179 => x"02bfccf1",
  1180 => x"f1c287cb",
  1181 => x"c648bfd0",
  1182 => x"d4f1c280",
  1183 => x"c4497358",
  1184 => x"264b2687",
  1185 => x"5b5e0e4f",
  1186 => x"f00e5d5c",
  1187 => x"59a6d086",
  1188 => x"4df4e3c2",
  1189 => x"f1c24cc0",
  1190 => x"78c148cc",
  1191 => x"c048a6c4",
  1192 => x"c27e7578",
  1193 => x"48bfd0f1",
  1194 => x"c006a8c0",
  1195 => x"7e7587fa",
  1196 => x"48f4e3c2",
  1197 => x"efc00298",
  1198 => x"c1fbc087",
  1199 => x"0266c81e",
  1200 => x"4dc087c4",
  1201 => x"4dc187c2",
  1202 => x"c9e44975",
  1203 => x"7086c487",
  1204 => x"c484c17e",
  1205 => x"80c14866",
  1206 => x"c258a6c8",
  1207 => x"acbfd0f1",
  1208 => x"6e87c503",
  1209 => x"87d1ff05",
  1210 => x"4cc04d6e",
  1211 => x"c3029d75",
  1212 => x"fbc087de",
  1213 => x"66c81ec1",
  1214 => x"cc87c702",
  1215 => x"78c048a6",
  1216 => x"a6cc87c5",
  1217 => x"cc78c148",
  1218 => x"c9e34966",
  1219 => x"7086c487",
  1220 => x"0298487e",
  1221 => x"4987e6c2",
  1222 => x"699781cb",
  1223 => x"0299d049",
  1224 => x"c187d6c1",
  1225 => x"744ae7c7",
  1226 => x"c191cc49",
  1227 => x"7281e8ec",
  1228 => x"c381c879",
  1229 => x"497451ff",
  1230 => x"f1c291de",
  1231 => x"85714de0",
  1232 => x"7d97c1c2",
  1233 => x"c049a5c1",
  1234 => x"ecc251e0",
  1235 => x"02bf97c4",
  1236 => x"84c187d2",
  1237 => x"c24ba5c2",
  1238 => x"db4ac4ec",
  1239 => x"c3f7fe49",
  1240 => x"87d9c187",
  1241 => x"c049a5cd",
  1242 => x"c284c151",
  1243 => x"4a6e4ba5",
  1244 => x"f6fe49cb",
  1245 => x"c4c187ee",
  1246 => x"cc497487",
  1247 => x"e8ecc191",
  1248 => x"dac5c181",
  1249 => x"c4ecc279",
  1250 => x"d802bf97",
  1251 => x"de497487",
  1252 => x"c284c191",
  1253 => x"714be0f1",
  1254 => x"c4ecc283",
  1255 => x"fe49dd4a",
  1256 => x"d887c1f6",
  1257 => x"de4b7487",
  1258 => x"e0f1c293",
  1259 => x"49a3cb83",
  1260 => x"84c151c0",
  1261 => x"cb4a6e73",
  1262 => x"e7f5fe49",
  1263 => x"4866c487",
  1264 => x"a6c880c1",
  1265 => x"03acc758",
  1266 => x"6e87c5c0",
  1267 => x"87e2fc05",
  1268 => x"c003acc7",
  1269 => x"f1c287e6",
  1270 => x"78c048cc",
  1271 => x"4adac5c1",
  1272 => x"91cc4974",
  1273 => x"81e8ecc1",
  1274 => x"49747972",
  1275 => x"f1c291de",
  1276 => x"51c081e0",
  1277 => x"acc784c1",
  1278 => x"87daff04",
  1279 => x"48c4eec1",
  1280 => x"80f750c0",
  1281 => x"40f1d1c1",
  1282 => x"78e4d0c1",
  1283 => x"c8c180c8",
  1284 => x"66cc78cf",
  1285 => x"e3fac049",
  1286 => x"268ef087",
  1287 => x"264c264d",
  1288 => x"004f264b",
  1289 => x"61422080",
  1290 => x"1e006b63",
  1291 => x"4b711e73",
  1292 => x"c191cc49",
  1293 => x"c881e8ec",
  1294 => x"ecc14aa1",
  1295 => x"501248dc",
  1296 => x"c04aa1c9",
  1297 => x"1248e0fd",
  1298 => x"c181ca50",
  1299 => x"1148e0ec",
  1300 => x"e0ecc150",
  1301 => x"1e49bf97",
  1302 => x"faf249c0",
  1303 => x"f8497387",
  1304 => x"8efc87e3",
  1305 => x"4f264b26",
  1306 => x"c049c01e",
  1307 => x"2687eefa",
  1308 => x"4a711e4f",
  1309 => x"c191cc49",
  1310 => x"c881e8ec",
  1311 => x"ecf0c281",
  1312 => x"c0501148",
  1313 => x"fe49a2f0",
  1314 => x"c087c1f0",
  1315 => x"87c7d749",
  1316 => x"ff1e4f26",
  1317 => x"ffc34ad4",
  1318 => x"48d0ff7a",
  1319 => x"de78e1c0",
  1320 => x"487a717a",
  1321 => x"7028b7c8",
  1322 => x"d048717a",
  1323 => x"7a7028b7",
  1324 => x"b7d84871",
  1325 => x"ff7a7028",
  1326 => x"e0c048d0",
  1327 => x"0e4f2678",
  1328 => x"5d5c5b5e",
  1329 => x"7186f40e",
  1330 => x"91cc494d",
  1331 => x"81e8ecc1",
  1332 => x"ca4aa1c8",
  1333 => x"a6c47ea1",
  1334 => x"e8f0c248",
  1335 => x"976e78bf",
  1336 => x"66c44bbf",
  1337 => x"122c734c",
  1338 => x"58a6cc48",
  1339 => x"84c19c70",
  1340 => x"699781c9",
  1341 => x"04acb749",
  1342 => x"4cc087c2",
  1343 => x"4abf976e",
  1344 => x"724966c8",
  1345 => x"c4b9ff31",
  1346 => x"48749966",
  1347 => x"4a703072",
  1348 => x"ecf0c2b1",
  1349 => x"f9fd7159",
  1350 => x"c21ec787",
  1351 => x"1ebfc8f1",
  1352 => x"1ee8ecc1",
  1353 => x"97ecf0c2",
  1354 => x"f4c149bf",
  1355 => x"c0497587",
  1356 => x"e887c9f6",
  1357 => x"264d268e",
  1358 => x"264b264c",
  1359 => x"1e731e4f",
  1360 => x"fd494b71",
  1361 => x"497387f9",
  1362 => x"2687f4fd",
  1363 => x"1e4f264b",
  1364 => x"4b711e73",
  1365 => x"024aa3c2",
  1366 => x"8ac187d6",
  1367 => x"87e2c005",
  1368 => x"bfc8f1c2",
  1369 => x"4887db02",
  1370 => x"f1c288c1",
  1371 => x"87d258cc",
  1372 => x"bfccf1c2",
  1373 => x"c287cb02",
  1374 => x"48bfc8f1",
  1375 => x"f1c280c1",
  1376 => x"1ec758cc",
  1377 => x"bfc8f1c2",
  1378 => x"e8ecc11e",
  1379 => x"ecf0c21e",
  1380 => x"cc49bf97",
  1381 => x"c0497387",
  1382 => x"f487e1f4",
  1383 => x"264b268e",
  1384 => x"5b5e0e4f",
  1385 => x"ff0e5d5c",
  1386 => x"e4c086cc",
  1387 => x"a6cc59a6",
  1388 => x"c478c048",
  1389 => x"c478c080",
  1390 => x"66c8c180",
  1391 => x"c180c478",
  1392 => x"c180c478",
  1393 => x"ccf1c278",
  1394 => x"e078c148",
  1395 => x"c8e187ee",
  1396 => x"87dde087",
  1397 => x"fbc04c70",
  1398 => x"f3c102ac",
  1399 => x"66e0c087",
  1400 => x"87e8c105",
  1401 => x"4a66c4c1",
  1402 => x"7e6a82c4",
  1403 => x"48f8e8c1",
  1404 => x"4120496e",
  1405 => x"51104120",
  1406 => x"4866c4c1",
  1407 => x"78ebd0c1",
  1408 => x"81c7496a",
  1409 => x"c4c15174",
  1410 => x"81c84966",
  1411 => x"a6d851c1",
  1412 => x"c178c248",
  1413 => x"c94966c4",
  1414 => x"c151c081",
  1415 => x"ca4966c4",
  1416 => x"c151c081",
  1417 => x"6a1ed81e",
  1418 => x"ff81c849",
  1419 => x"c887fedf",
  1420 => x"66c8c186",
  1421 => x"01a8c048",
  1422 => x"a6d087c7",
  1423 => x"cf78c148",
  1424 => x"66c8c187",
  1425 => x"d888c148",
  1426 => x"87c458a6",
  1427 => x"87c9dfff",
  1428 => x"cd029c74",
  1429 => x"66d087d9",
  1430 => x"66ccc148",
  1431 => x"cecd03a8",
  1432 => x"48a6c887",
  1433 => x"ff7e78c0",
  1434 => x"7087c6de",
  1435 => x"acd0c14c",
  1436 => x"87e7c205",
  1437 => x"6e48a6c4",
  1438 => x"87dce078",
  1439 => x"cc487e70",
  1440 => x"c506a866",
  1441 => x"48a6cc87",
  1442 => x"ddff786e",
  1443 => x"4c7087e3",
  1444 => x"05acecc0",
  1445 => x"d087eec1",
  1446 => x"91cc4966",
  1447 => x"8166c4c1",
  1448 => x"6a4aa1c4",
  1449 => x"4aa1c84d",
  1450 => x"d1c1526e",
  1451 => x"dcff79f1",
  1452 => x"4c7087ff",
  1453 => x"87d9029c",
  1454 => x"02acfbc0",
  1455 => x"557487d3",
  1456 => x"87eddcff",
  1457 => x"029c4c70",
  1458 => x"fbc087c7",
  1459 => x"edff05ac",
  1460 => x"55e0c087",
  1461 => x"c055c1c2",
  1462 => x"e0c07d97",
  1463 => x"66c44866",
  1464 => x"87db05a8",
  1465 => x"d44866d0",
  1466 => x"ca04a866",
  1467 => x"4866d087",
  1468 => x"a6d480c1",
  1469 => x"d487c858",
  1470 => x"88c14866",
  1471 => x"ff58a6d8",
  1472 => x"7087eedb",
  1473 => x"acd0c14c",
  1474 => x"dc87c905",
  1475 => x"80c14866",
  1476 => x"58a6e0c0",
  1477 => x"02acd0c1",
  1478 => x"6e87d9fd",
  1479 => x"66e0c048",
  1480 => x"eac905a8",
  1481 => x"a6e4c087",
  1482 => x"7478c048",
  1483 => x"88fbc048",
  1484 => x"7058a6c8",
  1485 => x"dcc90298",
  1486 => x"88cb4887",
  1487 => x"7058a6c8",
  1488 => x"cec10298",
  1489 => x"88c94887",
  1490 => x"7058a6c8",
  1491 => x"fec30298",
  1492 => x"88c44887",
  1493 => x"7058a6c8",
  1494 => x"87cf0298",
  1495 => x"c888c148",
  1496 => x"987058a6",
  1497 => x"87e7c302",
  1498 => x"c887dbc8",
  1499 => x"f0c048a6",
  1500 => x"fcd9ff78",
  1501 => x"c04c7087",
  1502 => x"c302acec",
  1503 => x"5ca6cc87",
  1504 => x"02acecc0",
  1505 => x"d9ff87cd",
  1506 => x"4c7087e7",
  1507 => x"05acecc0",
  1508 => x"c087f3ff",
  1509 => x"c002acec",
  1510 => x"d9ff87c4",
  1511 => x"1ec087d3",
  1512 => x"66d81eca",
  1513 => x"c191cc49",
  1514 => x"714866cc",
  1515 => x"58a6cc80",
  1516 => x"c44866c8",
  1517 => x"58a6d080",
  1518 => x"49bf66cc",
  1519 => x"87edd9ff",
  1520 => x"1ede1ec1",
  1521 => x"49bf66d4",
  1522 => x"87e1d9ff",
  1523 => x"497086d0",
  1524 => x"8808c048",
  1525 => x"58a6ecc0",
  1526 => x"c006a8c0",
  1527 => x"e8c087ee",
  1528 => x"a8dd4866",
  1529 => x"87e4c003",
  1530 => x"49bf66c4",
  1531 => x"8166e8c0",
  1532 => x"c051e0c0",
  1533 => x"c14966e8",
  1534 => x"bf66c481",
  1535 => x"51c1c281",
  1536 => x"4966e8c0",
  1537 => x"66c481c2",
  1538 => x"51c081bf",
  1539 => x"d0c1486e",
  1540 => x"496e78eb",
  1541 => x"66d881c8",
  1542 => x"c9496e51",
  1543 => x"5166dc81",
  1544 => x"81ca496e",
  1545 => x"d85166c8",
  1546 => x"80c14866",
  1547 => x"d058a6dc",
  1548 => x"66d44866",
  1549 => x"cbc004a8",
  1550 => x"4866d087",
  1551 => x"a6d480c1",
  1552 => x"87d1c558",
  1553 => x"c14866d4",
  1554 => x"58a6d888",
  1555 => x"ff87c6c5",
  1556 => x"c087c5d9",
  1557 => x"ff58a6ec",
  1558 => x"c087fdd8",
  1559 => x"c058a6f0",
  1560 => x"c005a8ec",
  1561 => x"48a687c9",
  1562 => x"7866e8c0",
  1563 => x"ff87c4c0",
  1564 => x"d087fed5",
  1565 => x"91cc4966",
  1566 => x"4866c4c1",
  1567 => x"a6c88071",
  1568 => x"4a66c458",
  1569 => x"66c482c8",
  1570 => x"c081ca49",
  1571 => x"c05166e8",
  1572 => x"c14966ec",
  1573 => x"66e8c081",
  1574 => x"7148c189",
  1575 => x"c1497030",
  1576 => x"7a977189",
  1577 => x"bfe8f0c2",
  1578 => x"66e8c049",
  1579 => x"4a6a9729",
  1580 => x"c0987148",
  1581 => x"c458a6f4",
  1582 => x"80c44866",
  1583 => x"c858a6cc",
  1584 => x"c04dbf66",
  1585 => x"6e4866e0",
  1586 => x"c5c002a8",
  1587 => x"c07ec087",
  1588 => x"7ec187c2",
  1589 => x"e0c01e6e",
  1590 => x"ff49751e",
  1591 => x"c887ced5",
  1592 => x"c04c7086",
  1593 => x"c106acb7",
  1594 => x"857487d4",
  1595 => x"49bf66c8",
  1596 => x"7581e0c0",
  1597 => x"e9c14b89",
  1598 => x"fe714ac4",
  1599 => x"c287e5e0",
  1600 => x"c07e7585",
  1601 => x"c14866e4",
  1602 => x"a6e8c080",
  1603 => x"66f0c058",
  1604 => x"7081c149",
  1605 => x"c5c002a9",
  1606 => x"c04dc087",
  1607 => x"4dc187c2",
  1608 => x"66cc1e75",
  1609 => x"e0c049bf",
  1610 => x"8966c481",
  1611 => x"66c81e71",
  1612 => x"f8d3ff49",
  1613 => x"c086c887",
  1614 => x"ff01a8b7",
  1615 => x"e4c087c5",
  1616 => x"d3c00266",
  1617 => x"4966c487",
  1618 => x"e4c081c9",
  1619 => x"66c45166",
  1620 => x"ffd2c148",
  1621 => x"87cec078",
  1622 => x"c94966c4",
  1623 => x"c451c281",
  1624 => x"d4c14866",
  1625 => x"66d078fd",
  1626 => x"a866d448",
  1627 => x"87cbc004",
  1628 => x"c14866d0",
  1629 => x"58a6d480",
  1630 => x"d487dac0",
  1631 => x"88c14866",
  1632 => x"c058a6d8",
  1633 => x"d2ff87cf",
  1634 => x"4c7087cf",
  1635 => x"ff87c6c0",
  1636 => x"7087c6d2",
  1637 => x"4866dc4c",
  1638 => x"e0c080c1",
  1639 => x"9c7458a6",
  1640 => x"87cbc002",
  1641 => x"c14866d0",
  1642 => x"04a866cc",
  1643 => x"d087f2f2",
  1644 => x"a8c74866",
  1645 => x"87e1c003",
  1646 => x"c24c66d0",
  1647 => x"c048ccf1",
  1648 => x"cc497478",
  1649 => x"66c4c191",
  1650 => x"4aa1c481",
  1651 => x"52c04a6a",
  1652 => x"c784c179",
  1653 => x"e2ff04ac",
  1654 => x"66e0c087",
  1655 => x"87e2c002",
  1656 => x"4966c4c1",
  1657 => x"c181d4c1",
  1658 => x"c14a66c4",
  1659 => x"52c082dc",
  1660 => x"79f1d1c1",
  1661 => x"4966c4c1",
  1662 => x"c181d8c1",
  1663 => x"c079c8e9",
  1664 => x"c4c187d6",
  1665 => x"d4c14966",
  1666 => x"66c4c181",
  1667 => x"82d8c14a",
  1668 => x"7ad0e9c1",
  1669 => x"79e8d1c1",
  1670 => x"4966c4c1",
  1671 => x"c181e0c1",
  1672 => x"ff79cfd5",
  1673 => x"cc87e9cf",
  1674 => x"ccff4866",
  1675 => x"264d268e",
  1676 => x"264b264c",
  1677 => x"0000004f",
  1678 => x"64616f4c",
  1679 => x"202e2a20",
  1680 => x"00000000",
  1681 => x"0000203a",
  1682 => x"61422080",
  1683 => x"00006b63",
  1684 => x"78452080",
  1685 => x"1e007469",
  1686 => x"f1c21ec7",
  1687 => x"c11ebfc8",
  1688 => x"c21ee8ec",
  1689 => x"bf97ecf0",
  1690 => x"87f5ec49",
  1691 => x"49e8ecc1",
  1692 => x"87d6e2c0",
  1693 => x"4f268ef4",
  1694 => x"c81e731e",
  1695 => x"eec187c3",
  1696 => x"ecc148c0",
  1697 => x"e8fe78c8",
  1698 => x"e1c049a0",
  1699 => x"49c787fc",
  1700 => x"87e8e0c0",
  1701 => x"e2c049c1",
  1702 => x"d4ff87c3",
  1703 => x"78ffc348",
  1704 => x"48d4f1c2",
  1705 => x"e3fe50c0",
  1706 => x"987087e2",
  1707 => x"fe87cd02",
  1708 => x"7087deed",
  1709 => x"87c40298",
  1710 => x"87c24ac1",
  1711 => x"9a724ac0",
  1712 => x"c187c802",
  1713 => x"fe49d4ec",
  1714 => x"c287dcd7",
  1715 => x"c048c8f1",
  1716 => x"ecf0c278",
  1717 => x"4950c048",
  1718 => x"c087fcfd",
  1719 => x"7087cdf6",
  1720 => x"cb029b4b",
  1721 => x"c4eec187",
  1722 => x"df49c75b",
  1723 => x"87c687ce",
  1724 => x"e0c049c0",
  1725 => x"c2c387e7",
  1726 => x"c8e2c087",
  1727 => x"d4f0c087",
  1728 => x"87f5ff87",
  1729 => x"4f264b26",
  1730 => x"746f6f42",
  1731 => x"2e676e69",
  1732 => x"00002e2e",
  1733 => x"4f204453",
  1734 => x"0000004b",
  1735 => x"00000000",
  1736 => x"00000000",
  1737 => x"00000001",
  1738 => x"0000115a",
  1739 => x"00002c60",
  1740 => x"00000000",
  1741 => x"0000115a",
  1742 => x"00002c7e",
  1743 => x"00000000",
  1744 => x"0000115a",
  1745 => x"00002c9c",
  1746 => x"00000000",
  1747 => x"0000115a",
  1748 => x"00002cba",
  1749 => x"00000000",
  1750 => x"0000115a",
  1751 => x"00002cd8",
  1752 => x"00000000",
  1753 => x"0000115a",
  1754 => x"00002cf6",
  1755 => x"00000000",
  1756 => x"0000115a",
  1757 => x"00002d14",
  1758 => x"00000000",
  1759 => x"00001471",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"0000120f",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"db86fc1e",
  1766 => x"fc7e7087",
  1767 => x"1e4f268e",
  1768 => x"c048f0fe",
  1769 => x"7909cd78",
  1770 => x"1e4f2609",
  1771 => x"49d4eec1",
  1772 => x"4f2687ed",
  1773 => x"bff0fe1e",
  1774 => x"1e4f2648",
  1775 => x"c148f0fe",
  1776 => x"1e4f2678",
  1777 => x"c048f0fe",
  1778 => x"1e4f2678",
  1779 => x"52c04a71",
  1780 => x"0e4f2651",
  1781 => x"5d5c5b5e",
  1782 => x"7186f40e",
  1783 => x"7e6d974d",
  1784 => x"974ca5c1",
  1785 => x"a6c8486c",
  1786 => x"c4486e58",
  1787 => x"c505a866",
  1788 => x"c048ff87",
  1789 => x"caff87e6",
  1790 => x"49a5c287",
  1791 => x"714b6c97",
  1792 => x"6b974ba3",
  1793 => x"7e6c974b",
  1794 => x"80c1486e",
  1795 => x"c758a6c8",
  1796 => x"58a6cc98",
  1797 => x"fe7c9770",
  1798 => x"487387e1",
  1799 => x"4d268ef4",
  1800 => x"4b264c26",
  1801 => x"5e0e4f26",
  1802 => x"f40e5c5b",
  1803 => x"d84c7186",
  1804 => x"ffc34a66",
  1805 => x"4ba4c29a",
  1806 => x"73496c97",
  1807 => x"517249a1",
  1808 => x"6e7e6c97",
  1809 => x"c880c148",
  1810 => x"98c758a6",
  1811 => x"7058a6cc",
  1812 => x"268ef454",
  1813 => x"264b264c",
  1814 => x"86fc1e4f",
  1815 => x"e087e4fd",
  1816 => x"c0494abf",
  1817 => x"0299c0e0",
  1818 => x"1e7287cb",
  1819 => x"49f4f4c2",
  1820 => x"c487f3fe",
  1821 => x"87fcfc86",
  1822 => x"fefc7e70",
  1823 => x"268efc87",
  1824 => x"f4c21e4f",
  1825 => x"c2fd49f4",
  1826 => x"d9f1c187",
  1827 => x"87cffc49",
  1828 => x"2687edc3",
  1829 => x"5b5e0e4f",
  1830 => x"fc0e5d5c",
  1831 => x"ff7e7186",
  1832 => x"f4c24dd4",
  1833 => x"eafc49f4",
  1834 => x"c04b7087",
  1835 => x"c204abb7",
  1836 => x"f0c387f8",
  1837 => x"87c905ab",
  1838 => x"48f8f5c1",
  1839 => x"d9c278c1",
  1840 => x"abe0c387",
  1841 => x"c187c905",
  1842 => x"c148fcf5",
  1843 => x"87cac278",
  1844 => x"bffcf5c1",
  1845 => x"c287c602",
  1846 => x"c24ca3c0",
  1847 => x"c14c7387",
  1848 => x"02bff8f5",
  1849 => x"7487e0c0",
  1850 => x"29b7c449",
  1851 => x"d4f7c191",
  1852 => x"cf4a7481",
  1853 => x"c192c29a",
  1854 => x"70307248",
  1855 => x"72baff4a",
  1856 => x"70986948",
  1857 => x"7487db79",
  1858 => x"29b7c449",
  1859 => x"d4f7c191",
  1860 => x"cf4a7481",
  1861 => x"c392c29a",
  1862 => x"70307248",
  1863 => x"b069484a",
  1864 => x"056e7970",
  1865 => x"ff87e7c0",
  1866 => x"e1c848d0",
  1867 => x"c17dc578",
  1868 => x"02bffcf5",
  1869 => x"e0c387c3",
  1870 => x"f8f5c17d",
  1871 => x"87c302bf",
  1872 => x"737df0c3",
  1873 => x"48d0ff7d",
  1874 => x"c078e1c8",
  1875 => x"f5c178e0",
  1876 => x"78c048fc",
  1877 => x"48f8f5c1",
  1878 => x"f4c278c0",
  1879 => x"f2f949f4",
  1880 => x"c04b7087",
  1881 => x"fd03abb7",
  1882 => x"48c087c8",
  1883 => x"4d268efc",
  1884 => x"4b264c26",
  1885 => x"00004f26",
  1886 => x"00000000",
  1887 => x"00000000",
  1888 => x"724ac01e",
  1889 => x"c191c449",
  1890 => x"c081d4f7",
  1891 => x"d082c179",
  1892 => x"ee04aab7",
  1893 => x"0e4f2687",
  1894 => x"5d5c5b5e",
  1895 => x"f84d710e",
  1896 => x"4a7587e1",
  1897 => x"922ab7c4",
  1898 => x"82d4f7c1",
  1899 => x"9ccf4c75",
  1900 => x"496a94c2",
  1901 => x"c32b744b",
  1902 => x"7448c29b",
  1903 => x"ff4c7030",
  1904 => x"714874bc",
  1905 => x"f77a7098",
  1906 => x"487387f1",
  1907 => x"4c264d26",
  1908 => x"4f264b26",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"00000000",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"48d0ff1e",
  1926 => x"7178e1c8",
  1927 => x"08d4ff48",
  1928 => x"1e4f2678",
  1929 => x"c848d0ff",
  1930 => x"487178e1",
  1931 => x"7808d4ff",
  1932 => x"ff4866c4",
  1933 => x"267808d4",
  1934 => x"4a711e4f",
  1935 => x"1e4966c4",
  1936 => x"deff4972",
  1937 => x"48d0ff87",
  1938 => x"fc78e0c0",
  1939 => x"1e4f268e",
  1940 => x"4b711e73",
  1941 => x"1e4966c8",
  1942 => x"e0c14a73",
  1943 => x"d8ff49a2",
  1944 => x"268efc87",
  1945 => x"1e4f264b",
  1946 => x"c848d0ff",
  1947 => x"487178c9",
  1948 => x"7808d4ff",
  1949 => x"711e4f26",
  1950 => x"87eb494a",
  1951 => x"c848d0ff",
  1952 => x"1e4f2678",
  1953 => x"4b711e73",
  1954 => x"bfccf5c2",
  1955 => x"c287c302",
  1956 => x"d0ff87eb",
  1957 => x"78c9c848",
  1958 => x"e0c04873",
  1959 => x"08d4ffb0",
  1960 => x"c0f5c278",
  1961 => x"c878c048",
  1962 => x"87c50266",
  1963 => x"c249ffc3",
  1964 => x"c249c087",
  1965 => x"cc59c8f5",
  1966 => x"87c60266",
  1967 => x"4ad5d5c5",
  1968 => x"ffcf87c4",
  1969 => x"f5c24aff",
  1970 => x"f5c25acc",
  1971 => x"78c148cc",
  1972 => x"4f264b26",
  1973 => x"5c5b5e0e",
  1974 => x"4d710e5d",
  1975 => x"bfc8f5c2",
  1976 => x"029d754b",
  1977 => x"c84987cb",
  1978 => x"fcf9c191",
  1979 => x"c482714a",
  1980 => x"fcfdc187",
  1981 => x"124cc04a",
  1982 => x"c2997349",
  1983 => x"48bfc4f5",
  1984 => x"d4ffb871",
  1985 => x"b7c17808",
  1986 => x"b7c8842b",
  1987 => x"87e704ac",
  1988 => x"bfc0f5c2",
  1989 => x"c280c848",
  1990 => x"2658c4f5",
  1991 => x"264c264d",
  1992 => x"1e4f264b",
  1993 => x"4b711e73",
  1994 => x"029a4a13",
  1995 => x"497287cb",
  1996 => x"1387e1fe",
  1997 => x"f5059a4a",
  1998 => x"264b2687",
  1999 => x"f5c21e4f",
  2000 => x"c249bfc0",
  2001 => x"c148c0f5",
  2002 => x"c0c478a1",
  2003 => x"db03a9b7",
  2004 => x"48d4ff87",
  2005 => x"bfc4f5c2",
  2006 => x"c0f5c278",
  2007 => x"f5c249bf",
  2008 => x"a1c148c0",
  2009 => x"b7c0c478",
  2010 => x"87e504a9",
  2011 => x"c848d0ff",
  2012 => x"ccf5c278",
  2013 => x"2678c048",
  2014 => x"0000004f",
  2015 => x"00000000",
  2016 => x"00000000",
  2017 => x"5f000000",
  2018 => x"0000005f",
  2019 => x"00030300",
  2020 => x"00000303",
  2021 => x"147f7f14",
  2022 => x"00147f7f",
  2023 => x"6b2e2400",
  2024 => x"00123a6b",
  2025 => x"18366a4c",
  2026 => x"0032566c",
  2027 => x"594f7e30",
  2028 => x"40683a77",
  2029 => x"07040000",
  2030 => x"00000003",
  2031 => x"3e1c0000",
  2032 => x"00004163",
  2033 => x"63410000",
  2034 => x"00001c3e",
  2035 => x"1c3e2a08",
  2036 => x"082a3e1c",
  2037 => x"3e080800",
  2038 => x"0008083e",
  2039 => x"e0800000",
  2040 => x"00000060",
  2041 => x"08080800",
  2042 => x"00080808",
  2043 => x"60000000",
  2044 => x"00000060",
  2045 => x"18306040",
  2046 => x"0103060c",
  2047 => x"597f3e00",
  2048 => x"003e7f4d",
  2049 => x"7f060400",
  2050 => x"0000007f",
  2051 => x"71634200",
  2052 => x"00464f59",
  2053 => x"49632200",
  2054 => x"00367f49",
  2055 => x"13161c18",
  2056 => x"00107f7f",
  2057 => x"45672700",
  2058 => x"00397d45",
  2059 => x"4b7e3c00",
  2060 => x"00307949",
  2061 => x"71010100",
  2062 => x"00070f79",
  2063 => x"497f3600",
  2064 => x"00367f49",
  2065 => x"494f0600",
  2066 => x"001e3f69",
  2067 => x"66000000",
  2068 => x"00000066",
  2069 => x"e6800000",
  2070 => x"00000066",
  2071 => x"14080800",
  2072 => x"00222214",
  2073 => x"14141400",
  2074 => x"00141414",
  2075 => x"14222200",
  2076 => x"00080814",
  2077 => x"51030200",
  2078 => x"00060f59",
  2079 => x"5d417f3e",
  2080 => x"001e1f55",
  2081 => x"097f7e00",
  2082 => x"007e7f09",
  2083 => x"497f7f00",
  2084 => x"00367f49",
  2085 => x"633e1c00",
  2086 => x"00414141",
  2087 => x"417f7f00",
  2088 => x"001c3e63",
  2089 => x"497f7f00",
  2090 => x"00414149",
  2091 => x"097f7f00",
  2092 => x"00010109",
  2093 => x"417f3e00",
  2094 => x"007a7b49",
  2095 => x"087f7f00",
  2096 => x"007f7f08",
  2097 => x"7f410000",
  2098 => x"0000417f",
  2099 => x"40602000",
  2100 => x"003f7f40",
  2101 => x"1c087f7f",
  2102 => x"00416336",
  2103 => x"407f7f00",
  2104 => x"00404040",
  2105 => x"0c067f7f",
  2106 => x"007f7f06",
  2107 => x"0c067f7f",
  2108 => x"007f7f18",
  2109 => x"417f3e00",
  2110 => x"003e7f41",
  2111 => x"097f7f00",
  2112 => x"00060f09",
  2113 => x"61417f3e",
  2114 => x"00407e7f",
  2115 => x"097f7f00",
  2116 => x"00667f19",
  2117 => x"4d6f2600",
  2118 => x"00327b59",
  2119 => x"7f010100",
  2120 => x"0001017f",
  2121 => x"407f3f00",
  2122 => x"003f7f40",
  2123 => x"703f0f00",
  2124 => x"000f3f70",
  2125 => x"18307f7f",
  2126 => x"007f7f30",
  2127 => x"1c366341",
  2128 => x"4163361c",
  2129 => x"7c060301",
  2130 => x"0103067c",
  2131 => x"4d597161",
  2132 => x"00414347",
  2133 => x"7f7f0000",
  2134 => x"00004141",
  2135 => x"0c060301",
  2136 => x"40603018",
  2137 => x"41410000",
  2138 => x"00007f7f",
  2139 => x"03060c08",
  2140 => x"00080c06",
  2141 => x"80808080",
  2142 => x"00808080",
  2143 => x"03000000",
  2144 => x"00000407",
  2145 => x"54742000",
  2146 => x"00787c54",
  2147 => x"447f7f00",
  2148 => x"00387c44",
  2149 => x"447c3800",
  2150 => x"00004444",
  2151 => x"447c3800",
  2152 => x"007f7f44",
  2153 => x"547c3800",
  2154 => x"00185c54",
  2155 => x"7f7e0400",
  2156 => x"00000505",
  2157 => x"a4bc1800",
  2158 => x"007cfca4",
  2159 => x"047f7f00",
  2160 => x"00787c04",
  2161 => x"3d000000",
  2162 => x"0000407d",
  2163 => x"80808000",
  2164 => x"00007dfd",
  2165 => x"107f7f00",
  2166 => x"00446c38",
  2167 => x"3f000000",
  2168 => x"0000407f",
  2169 => x"180c7c7c",
  2170 => x"00787c0c",
  2171 => x"047c7c00",
  2172 => x"00787c04",
  2173 => x"447c3800",
  2174 => x"00387c44",
  2175 => x"24fcfc00",
  2176 => x"00183c24",
  2177 => x"243c1800",
  2178 => x"00fcfc24",
  2179 => x"047c7c00",
  2180 => x"00080c04",
  2181 => x"545c4800",
  2182 => x"00207454",
  2183 => x"7f3f0400",
  2184 => x"00004444",
  2185 => x"407c3c00",
  2186 => x"007c7c40",
  2187 => x"603c1c00",
  2188 => x"001c3c60",
  2189 => x"30607c3c",
  2190 => x"003c7c60",
  2191 => x"10386c44",
  2192 => x"00446c38",
  2193 => x"e0bc1c00",
  2194 => x"001c3c60",
  2195 => x"74644400",
  2196 => x"00444c5c",
  2197 => x"3e080800",
  2198 => x"00414177",
  2199 => x"7f000000",
  2200 => x"0000007f",
  2201 => x"77414100",
  2202 => x"0008083e",
  2203 => x"03010102",
  2204 => x"00010202",
  2205 => x"7f7f7f7f",
  2206 => x"007f7f7f",
  2207 => x"1c1c0808",
  2208 => x"7f7f3e3e",
  2209 => x"3e3e7f7f",
  2210 => x"08081c1c",
  2211 => x"7c181000",
  2212 => x"0010187c",
  2213 => x"7c301000",
  2214 => x"0010307c",
  2215 => x"60603010",
  2216 => x"00061e78",
  2217 => x"183c6642",
  2218 => x"0042663c",
  2219 => x"c26a3878",
  2220 => x"00386cc6",
  2221 => x"60000060",
  2222 => x"00600000",
  2223 => x"5c5b5e0e",
  2224 => x"86fc0e5d",
  2225 => x"f5c27e71",
  2226 => x"c04cbfd4",
  2227 => x"c41ec04b",
  2228 => x"c402ab66",
  2229 => x"c24dc087",
  2230 => x"754dc187",
  2231 => x"ee49731e",
  2232 => x"86c887e1",
  2233 => x"ef49e0c0",
  2234 => x"a4c487ea",
  2235 => x"f0496a4a",
  2236 => x"c8f187f1",
  2237 => x"c184cc87",
  2238 => x"abb7c883",
  2239 => x"87cdff04",
  2240 => x"4d268efc",
  2241 => x"4b264c26",
  2242 => x"711e4f26",
  2243 => x"d8f5c24a",
  2244 => x"d8f5c25a",
  2245 => x"4978c748",
  2246 => x"2687e1fe",
  2247 => x"1e731e4f",
  2248 => x"b7c04a71",
  2249 => x"87d303aa",
  2250 => x"bff8d9c2",
  2251 => x"c187c405",
  2252 => x"c087c24b",
  2253 => x"fcd9c24b",
  2254 => x"c287c45b",
  2255 => x"fc5afcd9",
  2256 => x"f8d9c248",
  2257 => x"c14a78bf",
  2258 => x"a2c0c19a",
  2259 => x"87e6ec49",
  2260 => x"4f264b26",
  2261 => x"c44a711e",
  2262 => x"49721e66",
  2263 => x"fc87f0eb",
  2264 => x"1e4f268e",
  2265 => x"c348d4ff",
  2266 => x"d0ff78ff",
  2267 => x"78e1c048",
  2268 => x"c148d4ff",
  2269 => x"c4487178",
  2270 => x"08d4ff30",
  2271 => x"48d0ff78",
  2272 => x"2678e0c0",
  2273 => x"5b5e0e4f",
  2274 => x"ec0e5d5c",
  2275 => x"48a6c886",
  2276 => x"c47e78c0",
  2277 => x"78bfec80",
  2278 => x"f5c280f8",
  2279 => x"e878bfd4",
  2280 => x"d9c24cbf",
  2281 => x"e349bff8",
  2282 => x"eecb87eb",
  2283 => x"87cccb49",
  2284 => x"c758a6d4",
  2285 => x"87dfe749",
  2286 => x"c9059870",
  2287 => x"4966cc87",
  2288 => x"c10299c1",
  2289 => x"66d087c4",
  2290 => x"ec7ec14d",
  2291 => x"d9c24bbf",
  2292 => x"e249bff8",
  2293 => x"497587ff",
  2294 => x"7087edca",
  2295 => x"87d70298",
  2296 => x"bfe0d9c2",
  2297 => x"c2b9c149",
  2298 => x"7159e4d9",
  2299 => x"cb87f4fd",
  2300 => x"c7ca49ee",
  2301 => x"c74d7087",
  2302 => x"87dbe649",
  2303 => x"ff059870",
  2304 => x"497387c7",
  2305 => x"fe0599c1",
  2306 => x"026e87ff",
  2307 => x"c287e3c0",
  2308 => x"4abff8d9",
  2309 => x"d9c2bac1",
  2310 => x"0afc5afc",
  2311 => x"9ac10a7a",
  2312 => x"49a2c0c1",
  2313 => x"c187cfe9",
  2314 => x"eae549da",
  2315 => x"48a6c887",
  2316 => x"d9c278c1",
  2317 => x"c105bff8",
  2318 => x"c0c887c5",
  2319 => x"d9c24dc0",
  2320 => x"49134be4",
  2321 => x"87cfe549",
  2322 => x"c2029870",
  2323 => x"c1b47587",
  2324 => x"ff052db7",
  2325 => x"497487ec",
  2326 => x"7199ffc3",
  2327 => x"fb49c01e",
  2328 => x"497487f2",
  2329 => x"7129b7c8",
  2330 => x"fb49c11e",
  2331 => x"86c887e6",
  2332 => x"e449fdc3",
  2333 => x"fac387e1",
  2334 => x"87dbe449",
  2335 => x"7487d4c7",
  2336 => x"99ffc349",
  2337 => x"712cb7c8",
  2338 => x"029c74b4",
  2339 => x"d9c287df",
  2340 => x"c749bff4",
  2341 => x"987087f2",
  2342 => x"87c4c005",
  2343 => x"87d34cc0",
  2344 => x"c749e0c2",
  2345 => x"d9c287d6",
  2346 => x"c6c058f8",
  2347 => x"f4d9c287",
  2348 => x"7478c048",
  2349 => x"0599c849",
  2350 => x"c387cec0",
  2351 => x"d6e349f5",
  2352 => x"c2497087",
  2353 => x"e7c00299",
  2354 => x"d8f5c287",
  2355 => x"cac002bf",
  2356 => x"88c14887",
  2357 => x"58dcf5c2",
  2358 => x"c487d0c0",
  2359 => x"e0c14a66",
  2360 => x"c0026a82",
  2361 => x"ff4b87c5",
  2362 => x"c80f7349",
  2363 => x"78c148a6",
  2364 => x"99c44974",
  2365 => x"87cec005",
  2366 => x"e249f2c3",
  2367 => x"497087d9",
  2368 => x"c00299c2",
  2369 => x"f5c287f0",
  2370 => x"487ebfd8",
  2371 => x"03a8b7c7",
  2372 => x"6e87cbc0",
  2373 => x"c280c148",
  2374 => x"c058dcf5",
  2375 => x"66c487d3",
  2376 => x"80e0c148",
  2377 => x"bf6e7e70",
  2378 => x"87c5c002",
  2379 => x"7349fe4b",
  2380 => x"48a6c80f",
  2381 => x"fdc378c1",
  2382 => x"87dbe149",
  2383 => x"99c24970",
  2384 => x"87e9c002",
  2385 => x"bfd8f5c2",
  2386 => x"87c9c002",
  2387 => x"48d8f5c2",
  2388 => x"d3c078c0",
  2389 => x"4866c487",
  2390 => x"7080e0c1",
  2391 => x"02bf6e7e",
  2392 => x"4b87c5c0",
  2393 => x"0f7349fd",
  2394 => x"c148a6c8",
  2395 => x"49fac378",
  2396 => x"7087e4e0",
  2397 => x"0299c249",
  2398 => x"c287edc0",
  2399 => x"48bfd8f5",
  2400 => x"03a8b7c7",
  2401 => x"c287c9c0",
  2402 => x"c748d8f5",
  2403 => x"87d3c078",
  2404 => x"c14866c4",
  2405 => x"7e7080e0",
  2406 => x"c002bf6e",
  2407 => x"fc4b87c5",
  2408 => x"c80f7349",
  2409 => x"78c148a6",
  2410 => x"f5c27ec0",
  2411 => x"50c048d0",
  2412 => x"c349eecb",
  2413 => x"a6d487c6",
  2414 => x"d0f5c258",
  2415 => x"c105bf97",
  2416 => x"497487de",
  2417 => x"0599f0c3",
  2418 => x"c187cdc0",
  2419 => x"dfff49da",
  2420 => x"987087c5",
  2421 => x"87c8c102",
  2422 => x"bfe87ec1",
  2423 => x"ffc3494b",
  2424 => x"2bb7c899",
  2425 => x"d9c2b371",
  2426 => x"ff49bff8",
  2427 => x"d087e6da",
  2428 => x"d3c24966",
  2429 => x"02987087",
  2430 => x"c287c6c0",
  2431 => x"c148d0f5",
  2432 => x"d0f5c250",
  2433 => x"c005bf97",
  2434 => x"497387d6",
  2435 => x"0599f0c3",
  2436 => x"c187c5ff",
  2437 => x"ddff49da",
  2438 => x"987087fd",
  2439 => x"87f8fe05",
  2440 => x"e0c0026e",
  2441 => x"48a6cc87",
  2442 => x"bfd8f5c2",
  2443 => x"4966cc78",
  2444 => x"66c491cc",
  2445 => x"70807148",
  2446 => x"02bf6e7e",
  2447 => x"4b87c6c0",
  2448 => x"734966cc",
  2449 => x"0266c80f",
  2450 => x"c287c8c0",
  2451 => x"49bfd8f5",
  2452 => x"ec87e9f1",
  2453 => x"264d268e",
  2454 => x"264b264c",
  2455 => x"0000004f",
  2456 => x"00000000",
  2457 => x"14111258",
  2458 => x"231c1b1d",
  2459 => x"9491595a",
  2460 => x"f4ebf2f5",
  2461 => x"00000000",
  2462 => x"00000000",
  2463 => x"ff4a711e",
  2464 => x"7249bfc8",
  2465 => x"4f2648a1",
  2466 => x"bfc8ff1e",
  2467 => x"c0c0fe89",
  2468 => x"a9c0c0c0",
  2469 => x"c087c401",
  2470 => x"c187c24a",
  2471 => x"2648724a",
  2472 => x"5b5e0e4f",
  2473 => x"710e5d5c",
  2474 => x"4cd4ff4b",
  2475 => x"c04866d0",
  2476 => x"ff49d678",
  2477 => x"c387dddd",
  2478 => x"496c7cff",
  2479 => x"7199ffc3",
  2480 => x"f0c3494d",
  2481 => x"a9e0c199",
  2482 => x"c387cb05",
  2483 => x"486c7cff",
  2484 => x"66d098c3",
  2485 => x"ffc37808",
  2486 => x"494a6c7c",
  2487 => x"ffc331c8",
  2488 => x"714a6c7c",
  2489 => x"c84972b2",
  2490 => x"7cffc331",
  2491 => x"b2714a6c",
  2492 => x"31c84972",
  2493 => x"6c7cffc3",
  2494 => x"ffb2714a",
  2495 => x"e0c048d0",
  2496 => x"029b7378",
  2497 => x"7b7287c2",
  2498 => x"4d264875",
  2499 => x"4b264c26",
  2500 => x"261e4f26",
  2501 => x"5b5e0e4f",
  2502 => x"86f80e5c",
  2503 => x"a6c81e76",
  2504 => x"87fdfd49",
  2505 => x"4b7086c4",
  2506 => x"a8c2486e",
  2507 => x"87f0c203",
  2508 => x"f0c34a73",
  2509 => x"aad0c19a",
  2510 => x"c187c702",
  2511 => x"c205aae0",
  2512 => x"497387de",
  2513 => x"c30299c8",
  2514 => x"87c6ff87",
  2515 => x"9cc34c73",
  2516 => x"c105acc2",
  2517 => x"66c487c2",
  2518 => x"7131c949",
  2519 => x"4a66c41e",
  2520 => x"f5c292d4",
  2521 => x"817249dc",
  2522 => x"87e8cdfe",
  2523 => x"daff49d8",
  2524 => x"c0c887e2",
  2525 => x"f4e3c21e",
  2526 => x"dae7fd49",
  2527 => x"48d0ff87",
  2528 => x"c278e0c0",
  2529 => x"cc1ef4e3",
  2530 => x"92d44a66",
  2531 => x"49dcf5c2",
  2532 => x"cbfe8172",
  2533 => x"86cc87ef",
  2534 => x"c105acc1",
  2535 => x"66c487c2",
  2536 => x"7131c949",
  2537 => x"4a66c41e",
  2538 => x"f5c292d4",
  2539 => x"817249dc",
  2540 => x"87e0ccfe",
  2541 => x"1ef4e3c2",
  2542 => x"d44a66c8",
  2543 => x"dcf5c292",
  2544 => x"fe817249",
  2545 => x"d787efc9",
  2546 => x"c7d9ff49",
  2547 => x"1ec0c887",
  2548 => x"49f4e3c2",
  2549 => x"87dce5fd",
  2550 => x"d0ff86cc",
  2551 => x"78e0c048",
  2552 => x"4c268ef8",
  2553 => x"4f264b26",
  2554 => x"5c5b5e0e",
  2555 => x"86fc0e5d",
  2556 => x"d4ff4d71",
  2557 => x"7e66d44c",
  2558 => x"a8b7c348",
  2559 => x"87e2c101",
  2560 => x"66c41e75",
  2561 => x"c293d44b",
  2562 => x"7383dcf5",
  2563 => x"e4c3fe49",
  2564 => x"49a3c887",
  2565 => x"d0ff4969",
  2566 => x"78e1c848",
  2567 => x"48717cdd",
  2568 => x"7098ffc3",
  2569 => x"c84a717c",
  2570 => x"48722ab7",
  2571 => x"7098ffc3",
  2572 => x"d04a717c",
  2573 => x"48722ab7",
  2574 => x"7098ffc3",
  2575 => x"d848717c",
  2576 => x"7c7028b7",
  2577 => x"7c7c7cc0",
  2578 => x"7c7c7c7c",
  2579 => x"7c7c7c7c",
  2580 => x"48d0ff7c",
  2581 => x"c478e0c0",
  2582 => x"49dc1e66",
  2583 => x"87d9d7ff",
  2584 => x"8efc86c8",
  2585 => x"4c264d26",
  2586 => x"4f264b26",
  2587 => x"c01e731e",
  2588 => x"e2c21e4b",
  2589 => x"fd49bfe8",
  2590 => x"86c487ee",
  2591 => x"bfece2c2",
  2592 => x"c1dcfe49",
  2593 => x"05987087",
  2594 => x"e2c287c4",
  2595 => x"48734bd4",
  2596 => x"4f264b26",
  2597 => x"204d4f52",
  2598 => x"64616f6c",
  2599 => x"20676e69",
  2600 => x"6c696166",
  2601 => x"00006465",
  2602 => x"000028b0",
  2603 => x"000028bc",
  2604 => x"20434242",
  2605 => x"20202020",
  2606 => x"00444856",
  2607 => x"20434242",
  2608 => x"20202020",
  2609 => x"004d4f52",
  2610 => x"00001bab",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
