
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"64",x"44",x"00",x"00"),
     1 => (x"44",x"4c",x"5c",x"74"),
     2 => (x"08",x"08",x"00",x"00"),
     3 => (x"41",x"41",x"77",x"3e"),
     4 => (x"00",x"00",x"00",x"00"),
     5 => (x"00",x"00",x"7f",x"7f"),
     6 => (x"41",x"41",x"00",x"00"),
     7 => (x"08",x"08",x"3e",x"77"),
     8 => (x"01",x"01",x"02",x"00"),
     9 => (x"01",x"02",x"02",x"03"),
    10 => (x"7f",x"7f",x"7f",x"00"),
    11 => (x"7f",x"7f",x"7f",x"7f"),
    12 => (x"1c",x"08",x"08",x"00"),
    13 => (x"7f",x"3e",x"3e",x"1c"),
    14 => (x"3e",x"7f",x"7f",x"7f"),
    15 => (x"08",x"1c",x"1c",x"3e"),
    16 => (x"18",x"10",x"00",x"08"),
    17 => (x"10",x"18",x"7c",x"7c"),
    18 => (x"30",x"10",x"00",x"00"),
    19 => (x"10",x"30",x"7c",x"7c"),
    20 => (x"60",x"30",x"10",x"00"),
    21 => (x"06",x"1e",x"78",x"60"),
    22 => (x"3c",x"66",x"42",x"00"),
    23 => (x"42",x"66",x"3c",x"18"),
    24 => (x"6a",x"38",x"78",x"00"),
    25 => (x"38",x"6c",x"c6",x"c2"),
    26 => (x"00",x"00",x"60",x"00"),
    27 => (x"60",x"00",x"00",x"60"),
    28 => (x"5b",x"5e",x"0e",x"00"),
    29 => (x"1e",x"0e",x"5d",x"5c"),
    30 => (x"ee",x"c2",x"4c",x"71"),
    31 => (x"c0",x"4d",x"bf",x"dd"),
    32 => (x"74",x"1e",x"c0",x"4b"),
    33 => (x"87",x"c7",x"02",x"ab"),
    34 => (x"c0",x"48",x"a6",x"c4"),
    35 => (x"c4",x"87",x"c5",x"78"),
    36 => (x"78",x"c1",x"48",x"a6"),
    37 => (x"73",x"1e",x"66",x"c4"),
    38 => (x"87",x"df",x"ee",x"49"),
    39 => (x"e0",x"c0",x"86",x"c8"),
    40 => (x"87",x"ee",x"ef",x"49"),
    41 => (x"6a",x"4a",x"a5",x"c4"),
    42 => (x"87",x"f0",x"f0",x"49"),
    43 => (x"cb",x"87",x"c6",x"f1"),
    44 => (x"c8",x"83",x"c1",x"85"),
    45 => (x"ff",x"04",x"ab",x"b7"),
    46 => (x"26",x"26",x"87",x"c7"),
    47 => (x"26",x"4c",x"26",x"4d"),
    48 => (x"1e",x"4f",x"26",x"4b"),
    49 => (x"ee",x"c2",x"4a",x"71"),
    50 => (x"ee",x"c2",x"5a",x"e1"),
    51 => (x"78",x"c7",x"48",x"e1"),
    52 => (x"87",x"dd",x"fe",x"49"),
    53 => (x"73",x"1e",x"4f",x"26"),
    54 => (x"c0",x"4a",x"71",x"1e"),
    55 => (x"d3",x"03",x"aa",x"b7"),
    56 => (x"d8",x"d3",x"c2",x"87"),
    57 => (x"87",x"c4",x"05",x"bf"),
    58 => (x"87",x"c2",x"4b",x"c1"),
    59 => (x"d3",x"c2",x"4b",x"c0"),
    60 => (x"87",x"c4",x"5b",x"dc"),
    61 => (x"5a",x"dc",x"d3",x"c2"),
    62 => (x"bf",x"d8",x"d3",x"c2"),
    63 => (x"c1",x"9a",x"c1",x"4a"),
    64 => (x"ec",x"49",x"a2",x"c0"),
    65 => (x"48",x"fc",x"87",x"e8"),
    66 => (x"bf",x"d8",x"d3",x"c2"),
    67 => (x"87",x"ef",x"fe",x"78"),
    68 => (x"c4",x"4a",x"71",x"1e"),
    69 => (x"49",x"72",x"1e",x"66"),
    70 => (x"26",x"87",x"f9",x"ea"),
    71 => (x"ff",x"1e",x"4f",x"26"),
    72 => (x"ff",x"c3",x"48",x"d4"),
    73 => (x"48",x"d0",x"ff",x"78"),
    74 => (x"ff",x"78",x"e1",x"c0"),
    75 => (x"78",x"c1",x"48",x"d4"),
    76 => (x"30",x"c4",x"48",x"71"),
    77 => (x"78",x"08",x"d4",x"ff"),
    78 => (x"c0",x"48",x"d0",x"ff"),
    79 => (x"4f",x"26",x"78",x"e0"),
    80 => (x"5c",x"5b",x"5e",x"0e"),
    81 => (x"86",x"f4",x"0e",x"5d"),
    82 => (x"c0",x"48",x"a6",x"c4"),
    83 => (x"bf",x"ec",x"4b",x"78"),
    84 => (x"dd",x"ee",x"c2",x"7e"),
    85 => (x"bf",x"e8",x"4d",x"bf"),
    86 => (x"d8",x"d3",x"c2",x"4c"),
    87 => (x"fe",x"e2",x"49",x"bf"),
    88 => (x"49",x"ee",x"cb",x"87"),
    89 => (x"cc",x"87",x"f9",x"cd"),
    90 => (x"49",x"c7",x"58",x"a6"),
    91 => (x"70",x"87",x"f3",x"e6"),
    92 => (x"87",x"c8",x"05",x"98"),
    93 => (x"99",x"c1",x"49",x"6e"),
    94 => (x"87",x"c3",x"c1",x"02"),
    95 => (x"bf",x"ec",x"4b",x"c1"),
    96 => (x"d8",x"d3",x"c2",x"7e"),
    97 => (x"d6",x"e2",x"49",x"bf"),
    98 => (x"49",x"66",x"c8",x"87"),
    99 => (x"70",x"87",x"dd",x"cd"),
   100 => (x"87",x"d8",x"02",x"98"),
   101 => (x"bf",x"c0",x"d3",x"c2"),
   102 => (x"c2",x"b9",x"c1",x"49"),
   103 => (x"71",x"59",x"c4",x"d3"),
   104 => (x"cb",x"87",x"fb",x"fd"),
   105 => (x"f7",x"cc",x"49",x"ee"),
   106 => (x"58",x"a6",x"cc",x"87"),
   107 => (x"f1",x"e5",x"49",x"c7"),
   108 => (x"05",x"98",x"70",x"87"),
   109 => (x"6e",x"87",x"c5",x"ff"),
   110 => (x"05",x"99",x"c1",x"49"),
   111 => (x"73",x"87",x"fd",x"fe"),
   112 => (x"87",x"d0",x"02",x"9b"),
   113 => (x"cd",x"fc",x"49",x"ff"),
   114 => (x"49",x"da",x"c1",x"87"),
   115 => (x"c4",x"87",x"d3",x"e5"),
   116 => (x"78",x"c1",x"48",x"a6"),
   117 => (x"bf",x"d8",x"d3",x"c2"),
   118 => (x"87",x"d9",x"c1",x"05"),
   119 => (x"c8",x"48",x"a6",x"c4"),
   120 => (x"c2",x"78",x"c0",x"c0"),
   121 => (x"6e",x"7e",x"c4",x"d3"),
   122 => (x"6e",x"49",x"bf",x"97"),
   123 => (x"70",x"80",x"c1",x"48"),
   124 => (x"ed",x"e4",x"71",x"7e"),
   125 => (x"02",x"98",x"70",x"87"),
   126 => (x"66",x"c4",x"87",x"c3"),
   127 => (x"48",x"66",x"c4",x"b4"),
   128 => (x"c8",x"28",x"b7",x"c1"),
   129 => (x"98",x"70",x"58",x"a6"),
   130 => (x"87",x"db",x"ff",x"05"),
   131 => (x"e4",x"49",x"fd",x"c3"),
   132 => (x"fa",x"c3",x"87",x"d0"),
   133 => (x"87",x"ca",x"e4",x"49"),
   134 => (x"ff",x"c3",x"49",x"74"),
   135 => (x"c0",x"1e",x"71",x"99"),
   136 => (x"87",x"ec",x"fb",x"49"),
   137 => (x"b7",x"c8",x"49",x"74"),
   138 => (x"c1",x"1e",x"71",x"29"),
   139 => (x"87",x"e0",x"fb",x"49"),
   140 => (x"f4",x"c8",x"86",x"c8"),
   141 => (x"c3",x"49",x"74",x"87"),
   142 => (x"b7",x"c8",x"99",x"ff"),
   143 => (x"74",x"b4",x"71",x"2c"),
   144 => (x"87",x"df",x"02",x"9c"),
   145 => (x"bf",x"d4",x"d3",x"c2"),
   146 => (x"87",x"e0",x"ca",x"49"),
   147 => (x"c0",x"05",x"98",x"70"),
   148 => (x"4c",x"c0",x"87",x"c4"),
   149 => (x"e0",x"c2",x"87",x"d3"),
   150 => (x"87",x"c4",x"ca",x"49"),
   151 => (x"58",x"d8",x"d3",x"c2"),
   152 => (x"c2",x"87",x"c6",x"c0"),
   153 => (x"c0",x"48",x"d4",x"d3"),
   154 => (x"c2",x"49",x"74",x"78"),
   155 => (x"ce",x"c0",x"05",x"99"),
   156 => (x"49",x"eb",x"c3",x"87"),
   157 => (x"70",x"87",x"eb",x"e2"),
   158 => (x"02",x"99",x"c2",x"49"),
   159 => (x"c1",x"87",x"cf",x"c0"),
   160 => (x"6e",x"7e",x"a5",x"d8"),
   161 => (x"c5",x"c0",x"02",x"bf"),
   162 => (x"49",x"fb",x"4b",x"87"),
   163 => (x"49",x"74",x"0f",x"73"),
   164 => (x"c0",x"05",x"99",x"c1"),
   165 => (x"f4",x"c3",x"87",x"ce"),
   166 => (x"87",x"c6",x"e2",x"49"),
   167 => (x"99",x"c2",x"49",x"70"),
   168 => (x"87",x"cf",x"c0",x"02"),
   169 => (x"7e",x"a5",x"d8",x"c1"),
   170 => (x"c0",x"02",x"bf",x"6e"),
   171 => (x"fa",x"4b",x"87",x"c5"),
   172 => (x"74",x"0f",x"73",x"49"),
   173 => (x"05",x"99",x"c8",x"49"),
   174 => (x"c3",x"87",x"ce",x"c0"),
   175 => (x"e1",x"e1",x"49",x"f5"),
   176 => (x"c2",x"49",x"70",x"87"),
   177 => (x"e5",x"c0",x"02",x"99"),
   178 => (x"e1",x"ee",x"c2",x"87"),
   179 => (x"ca",x"c0",x"02",x"bf"),
   180 => (x"88",x"c1",x"48",x"87"),
   181 => (x"58",x"e5",x"ee",x"c2"),
   182 => (x"c1",x"87",x"ce",x"c0"),
   183 => (x"6a",x"4a",x"a5",x"d8"),
   184 => (x"87",x"c5",x"c0",x"02"),
   185 => (x"73",x"49",x"ff",x"4b"),
   186 => (x"48",x"a6",x"c4",x"0f"),
   187 => (x"49",x"74",x"78",x"c1"),
   188 => (x"c0",x"05",x"99",x"c4"),
   189 => (x"f2",x"c3",x"87",x"ce"),
   190 => (x"87",x"e6",x"e0",x"49"),
   191 => (x"99",x"c2",x"49",x"70"),
   192 => (x"87",x"ec",x"c0",x"02"),
   193 => (x"bf",x"e1",x"ee",x"c2"),
   194 => (x"b7",x"c7",x"48",x"7e"),
   195 => (x"cb",x"c0",x"03",x"a8"),
   196 => (x"c1",x"48",x"6e",x"87"),
   197 => (x"e5",x"ee",x"c2",x"80"),
   198 => (x"87",x"cf",x"c0",x"58"),
   199 => (x"7e",x"a5",x"d8",x"c1"),
   200 => (x"c0",x"02",x"bf",x"6e"),
   201 => (x"fe",x"4b",x"87",x"c5"),
   202 => (x"c4",x"0f",x"73",x"49"),
   203 => (x"78",x"c1",x"48",x"a6"),
   204 => (x"ff",x"49",x"fd",x"c3"),
   205 => (x"70",x"87",x"eb",x"df"),
   206 => (x"02",x"99",x"c2",x"49"),
   207 => (x"c2",x"87",x"e5",x"c0"),
   208 => (x"02",x"bf",x"e1",x"ee"),
   209 => (x"c2",x"87",x"c9",x"c0"),
   210 => (x"c0",x"48",x"e1",x"ee"),
   211 => (x"87",x"cf",x"c0",x"78"),
   212 => (x"7e",x"a5",x"d8",x"c1"),
   213 => (x"c0",x"02",x"bf",x"6e"),
   214 => (x"fd",x"4b",x"87",x"c5"),
   215 => (x"c4",x"0f",x"73",x"49"),
   216 => (x"78",x"c1",x"48",x"a6"),
   217 => (x"ff",x"49",x"fa",x"c3"),
   218 => (x"70",x"87",x"f7",x"de"),
   219 => (x"02",x"99",x"c2",x"49"),
   220 => (x"c2",x"87",x"e9",x"c0"),
   221 => (x"48",x"bf",x"e1",x"ee"),
   222 => (x"03",x"a8",x"b7",x"c7"),
   223 => (x"c2",x"87",x"c9",x"c0"),
   224 => (x"c7",x"48",x"e1",x"ee"),
   225 => (x"87",x"cf",x"c0",x"78"),
   226 => (x"7e",x"a5",x"d8",x"c1"),
   227 => (x"c0",x"02",x"bf",x"6e"),
   228 => (x"fc",x"4b",x"87",x"c5"),
   229 => (x"c4",x"0f",x"73",x"49"),
   230 => (x"78",x"c1",x"48",x"a6"),
   231 => (x"ee",x"c2",x"4b",x"c0"),
   232 => (x"50",x"c0",x"48",x"dc"),
   233 => (x"c4",x"49",x"ee",x"cb"),
   234 => (x"a6",x"cc",x"87",x"f6"),
   235 => (x"dc",x"ee",x"c2",x"58"),
   236 => (x"c1",x"05",x"bf",x"97"),
   237 => (x"49",x"74",x"87",x"de"),
   238 => (x"05",x"99",x"f0",x"c3"),
   239 => (x"c1",x"87",x"cd",x"c0"),
   240 => (x"dd",x"ff",x"49",x"da"),
   241 => (x"98",x"70",x"87",x"dc"),
   242 => (x"87",x"c8",x"c1",x"02"),
   243 => (x"bf",x"e8",x"4b",x"c1"),
   244 => (x"ff",x"c3",x"49",x"4c"),
   245 => (x"2c",x"b7",x"c8",x"99"),
   246 => (x"d3",x"c2",x"b4",x"71"),
   247 => (x"ff",x"49",x"bf",x"d8"),
   248 => (x"c8",x"87",x"fc",x"d8"),
   249 => (x"c3",x"c4",x"49",x"66"),
   250 => (x"02",x"98",x"70",x"87"),
   251 => (x"c2",x"87",x"c6",x"c0"),
   252 => (x"c1",x"48",x"dc",x"ee"),
   253 => (x"dc",x"ee",x"c2",x"50"),
   254 => (x"c0",x"05",x"bf",x"97"),
   255 => (x"49",x"74",x"87",x"d6"),
   256 => (x"05",x"99",x"f0",x"c3"),
   257 => (x"c1",x"87",x"c5",x"ff"),
   258 => (x"dc",x"ff",x"49",x"da"),
   259 => (x"98",x"70",x"87",x"d4"),
   260 => (x"87",x"f8",x"fe",x"05"),
   261 => (x"c0",x"02",x"9b",x"73"),
   262 => (x"a6",x"c8",x"87",x"dc"),
   263 => (x"e1",x"ee",x"c2",x"48"),
   264 => (x"66",x"c8",x"78",x"bf"),
   265 => (x"75",x"91",x"cb",x"49"),
   266 => (x"bf",x"6e",x"7e",x"a1"),
   267 => (x"87",x"c6",x"c0",x"02"),
   268 => (x"49",x"66",x"c8",x"4b"),
   269 => (x"66",x"c4",x"0f",x"73"),
   270 => (x"87",x"c8",x"c0",x"02"),
   271 => (x"bf",x"e1",x"ee",x"c2"),
   272 => (x"87",x"ed",x"f0",x"49"),
   273 => (x"bf",x"dc",x"d3",x"c2"),
   274 => (x"87",x"dd",x"c0",x"02"),
   275 => (x"87",x"dc",x"c2",x"49"),
   276 => (x"c0",x"02",x"98",x"70"),
   277 => (x"ee",x"c2",x"87",x"d3"),
   278 => (x"f0",x"49",x"bf",x"e1"),
   279 => (x"49",x"c0",x"87",x"d3"),
   280 => (x"c2",x"87",x"f3",x"f1"),
   281 => (x"c0",x"48",x"dc",x"d3"),
   282 => (x"f1",x"8e",x"f4",x"78"),
   283 => (x"5e",x"0e",x"87",x"cd"),
   284 => (x"0e",x"5d",x"5c",x"5b"),
   285 => (x"c2",x"4c",x"71",x"1e"),
   286 => (x"49",x"bf",x"dd",x"ee"),
   287 => (x"4d",x"a1",x"cd",x"c1"),
   288 => (x"69",x"81",x"d1",x"c1"),
   289 => (x"02",x"9c",x"74",x"7e"),
   290 => (x"a5",x"c4",x"87",x"cf"),
   291 => (x"c2",x"7b",x"74",x"4b"),
   292 => (x"49",x"bf",x"dd",x"ee"),
   293 => (x"6e",x"87",x"ec",x"f0"),
   294 => (x"05",x"9c",x"74",x"7b"),
   295 => (x"4b",x"c0",x"87",x"c4"),
   296 => (x"4b",x"c1",x"87",x"c2"),
   297 => (x"ed",x"f0",x"49",x"73"),
   298 => (x"02",x"66",x"d4",x"87"),
   299 => (x"c0",x"49",x"87",x"c8"),
   300 => (x"4a",x"70",x"87",x"ee"),
   301 => (x"4a",x"c0",x"87",x"c2"),
   302 => (x"5a",x"e0",x"d3",x"c2"),
   303 => (x"87",x"fb",x"ef",x"26"),
   304 => (x"00",x"00",x"00",x"00"),
   305 => (x"14",x"11",x"12",x"58"),
   306 => (x"23",x"1c",x"1b",x"1d"),
   307 => (x"94",x"91",x"59",x"5a"),
   308 => (x"f4",x"eb",x"f2",x"f5"),
   309 => (x"00",x"00",x"00",x"00"),
   310 => (x"00",x"00",x"00",x"00"),
   311 => (x"00",x"00",x"00",x"00"),
   312 => (x"ff",x"4a",x"71",x"1e"),
   313 => (x"72",x"49",x"bf",x"c8"),
   314 => (x"4f",x"26",x"48",x"a1"),
   315 => (x"bf",x"c8",x"ff",x"1e"),
   316 => (x"c0",x"c0",x"fe",x"89"),
   317 => (x"a9",x"c0",x"c0",x"c0"),
   318 => (x"c0",x"87",x"c4",x"01"),
   319 => (x"c1",x"87",x"c2",x"4a"),
   320 => (x"26",x"48",x"72",x"4a"),
   321 => (x"5b",x"5e",x"0e",x"4f"),
   322 => (x"71",x"0e",x"5d",x"5c"),
   323 => (x"4c",x"d4",x"ff",x"4b"),
   324 => (x"c0",x"48",x"66",x"d0"),
   325 => (x"ff",x"49",x"d6",x"78"),
   326 => (x"c3",x"87",x"ff",x"d9"),
   327 => (x"49",x"6c",x"7c",x"ff"),
   328 => (x"71",x"99",x"ff",x"c3"),
   329 => (x"f0",x"c3",x"49",x"4d"),
   330 => (x"a9",x"e0",x"c1",x"99"),
   331 => (x"c3",x"87",x"cb",x"05"),
   332 => (x"48",x"6c",x"7c",x"ff"),
   333 => (x"66",x"d0",x"98",x"c3"),
   334 => (x"ff",x"c3",x"78",x"08"),
   335 => (x"49",x"4a",x"6c",x"7c"),
   336 => (x"ff",x"c3",x"31",x"c8"),
   337 => (x"71",x"4a",x"6c",x"7c"),
   338 => (x"c8",x"49",x"72",x"b2"),
   339 => (x"7c",x"ff",x"c3",x"31"),
   340 => (x"b2",x"71",x"4a",x"6c"),
   341 => (x"31",x"c8",x"49",x"72"),
   342 => (x"6c",x"7c",x"ff",x"c3"),
   343 => (x"ff",x"b2",x"71",x"4a"),
   344 => (x"e0",x"c0",x"48",x"d0"),
   345 => (x"02",x"9b",x"73",x"78"),
   346 => (x"7b",x"72",x"87",x"c2"),
   347 => (x"4d",x"26",x"48",x"75"),
   348 => (x"4b",x"26",x"4c",x"26"),
   349 => (x"26",x"1e",x"4f",x"26"),
   350 => (x"5b",x"5e",x"0e",x"4f"),
   351 => (x"86",x"f8",x"0e",x"5c"),
   352 => (x"a6",x"c8",x"1e",x"76"),
   353 => (x"87",x"fd",x"fd",x"49"),
   354 => (x"4b",x"70",x"86",x"c4"),
   355 => (x"a8",x"c2",x"48",x"6e"),
   356 => (x"87",x"f0",x"c2",x"03"),
   357 => (x"f0",x"c3",x"4a",x"73"),
   358 => (x"aa",x"d0",x"c1",x"9a"),
   359 => (x"c1",x"87",x"c7",x"02"),
   360 => (x"c2",x"05",x"aa",x"e0"),
   361 => (x"49",x"73",x"87",x"de"),
   362 => (x"c3",x"02",x"99",x"c8"),
   363 => (x"87",x"c6",x"ff",x"87"),
   364 => (x"9c",x"c3",x"4c",x"73"),
   365 => (x"c1",x"05",x"ac",x"c2"),
   366 => (x"66",x"c4",x"87",x"c2"),
   367 => (x"71",x"31",x"c9",x"49"),
   368 => (x"4a",x"66",x"c4",x"1e"),
   369 => (x"ee",x"c2",x"92",x"d4"),
   370 => (x"81",x"72",x"49",x"e5"),
   371 => (x"87",x"f7",x"cf",x"fe"),
   372 => (x"d7",x"ff",x"49",x"d8"),
   373 => (x"c0",x"c8",x"87",x"c4"),
   374 => (x"ce",x"dd",x"c2",x"1e"),
   375 => (x"fd",x"eb",x"fd",x"49"),
   376 => (x"48",x"d0",x"ff",x"87"),
   377 => (x"c2",x"78",x"e0",x"c0"),
   378 => (x"cc",x"1e",x"ce",x"dd"),
   379 => (x"92",x"d4",x"4a",x"66"),
   380 => (x"49",x"e5",x"ee",x"c2"),
   381 => (x"cd",x"fe",x"81",x"72"),
   382 => (x"86",x"cc",x"87",x"ff"),
   383 => (x"c1",x"05",x"ac",x"c1"),
   384 => (x"66",x"c4",x"87",x"c2"),
   385 => (x"71",x"31",x"c9",x"49"),
   386 => (x"4a",x"66",x"c4",x"1e"),
   387 => (x"ee",x"c2",x"92",x"d4"),
   388 => (x"81",x"72",x"49",x"e5"),
   389 => (x"87",x"ef",x"ce",x"fe"),
   390 => (x"1e",x"ce",x"dd",x"c2"),
   391 => (x"d4",x"4a",x"66",x"c8"),
   392 => (x"e5",x"ee",x"c2",x"92"),
   393 => (x"fe",x"81",x"72",x"49"),
   394 => (x"d7",x"87",x"c0",x"cc"),
   395 => (x"e9",x"d5",x"ff",x"49"),
   396 => (x"1e",x"c0",x"c8",x"87"),
   397 => (x"49",x"ce",x"dd",x"c2"),
   398 => (x"87",x"fb",x"e9",x"fd"),
   399 => (x"d0",x"ff",x"86",x"cc"),
   400 => (x"78",x"e0",x"c0",x"48"),
   401 => (x"e7",x"fc",x"8e",x"f8"),
   402 => (x"5b",x"5e",x"0e",x"87"),
   403 => (x"71",x"0e",x"5d",x"5c"),
   404 => (x"4c",x"d4",x"ff",x"4a"),
   405 => (x"c3",x"4d",x"66",x"d0"),
   406 => (x"c5",x"06",x"ad",x"b7"),
   407 => (x"c1",x"48",x"c0",x"87"),
   408 => (x"1e",x"72",x"87",x"e1"),
   409 => (x"93",x"d4",x"4b",x"75"),
   410 => (x"83",x"e5",x"ee",x"c2"),
   411 => (x"c6",x"fe",x"49",x"73"),
   412 => (x"83",x"c8",x"87",x"c7"),
   413 => (x"d0",x"ff",x"4b",x"6b"),
   414 => (x"78",x"e1",x"c8",x"48"),
   415 => (x"48",x"73",x"7c",x"dd"),
   416 => (x"70",x"98",x"ff",x"c3"),
   417 => (x"c8",x"49",x"73",x"7c"),
   418 => (x"48",x"71",x"29",x"b7"),
   419 => (x"70",x"98",x"ff",x"c3"),
   420 => (x"d0",x"49",x"73",x"7c"),
   421 => (x"48",x"71",x"29",x"b7"),
   422 => (x"70",x"98",x"ff",x"c3"),
   423 => (x"d8",x"48",x"73",x"7c"),
   424 => (x"7c",x"70",x"28",x"b7"),
   425 => (x"7c",x"7c",x"7c",x"c0"),
   426 => (x"7c",x"7c",x"7c",x"7c"),
   427 => (x"7c",x"7c",x"7c",x"7c"),
   428 => (x"48",x"d0",x"ff",x"7c"),
   429 => (x"75",x"78",x"e0",x"c0"),
   430 => (x"ff",x"49",x"dc",x"1e"),
   431 => (x"c8",x"87",x"c0",x"d4"),
   432 => (x"fa",x"48",x"73",x"86"),
   433 => (x"73",x"1e",x"87",x"e8"),
   434 => (x"1e",x"4b",x"c0",x"1e"),
   435 => (x"bf",x"c7",x"dc",x"c2"),
   436 => (x"87",x"f5",x"fd",x"49"),
   437 => (x"dc",x"c2",x"86",x"c4"),
   438 => (x"fe",x"49",x"bf",x"cb"),
   439 => (x"70",x"87",x"d0",x"dd"),
   440 => (x"87",x"c4",x"05",x"98"),
   441 => (x"4b",x"f4",x"db",x"c2"),
   442 => (x"87",x"c4",x"48",x"73"),
   443 => (x"4c",x"26",x"4d",x"26"),
   444 => (x"4f",x"26",x"4b",x"26"),
   445 => (x"20",x"4d",x"4f",x"52"),
   446 => (x"64",x"61",x"6f",x"6c"),
   447 => (x"20",x"67",x"6e",x"69"),
   448 => (x"6c",x"69",x"61",x"66"),
   449 => (x"0f",x"00",x"64",x"65"),
   450 => (x"1b",x"00",x"00",x"27"),
   451 => (x"42",x"00",x"00",x"27"),
   452 => (x"20",x"20",x"43",x"42"),
   453 => (x"56",x"20",x"20",x"20"),
   454 => (x"42",x"00",x"44",x"48"),
   455 => (x"20",x"20",x"43",x"42"),
   456 => (x"52",x"20",x"20",x"20"),
   457 => (x"52",x"00",x"4d",x"4f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

