library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c0f4c287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49c0f4c2",
    18 => x"48c8e1c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"c8e1c287",
    25 => x"c4e1c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e9c187f7",
    29 => x"e1c287c1",
    30 => x"e1c24dc8",
    31 => x"ad744cc8",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"731e741e",
    65 => x"c11e721e",
    66 => x"87d0048b",
    67 => x"02114812",
    68 => x"c34c87ca",
    69 => x"749c98df",
    70 => x"87eb0288",
    71 => x"4b264a26",
    72 => x"4f264c26",
    73 => x"8148731e",
    74 => x"c502a973",
    75 => x"05531287",
    76 => x"4f2687f6",
    77 => x"711e731e",
    78 => x"4b66c84a",
    79 => x"718bc149",
    80 => x"87cf0299",
    81 => x"d4ff4812",
    82 => x"49737808",
    83 => x"99718bc1",
    84 => x"2687f105",
    85 => x"0e4f264b",
    86 => x"0e5c5b5e",
    87 => x"d4ff4a71",
    88 => x"4b66cc4c",
    89 => x"718bc149",
    90 => x"87ce0299",
    91 => x"6c7cffc3",
    92 => x"c1497352",
    93 => x"0599718b",
    94 => x"4c2687f2",
    95 => x"4f264b26",
    96 => x"ff1e731e",
    97 => x"ffc34bd4",
    98 => x"c34a6b7b",
    99 => x"496b7bff",
   100 => x"b17232c8",
   101 => x"6b7bffc3",
   102 => x"7131c84a",
   103 => x"7bffc3b2",
   104 => x"32c8496b",
   105 => x"4871b172",
   106 => x"4f264b26",
   107 => x"5c5b5e0e",
   108 => x"4d710e5d",
   109 => x"754cd4ff",
   110 => x"98ffc348",
   111 => x"e1c27c70",
   112 => x"c805bfc8",
   113 => x"4866d087",
   114 => x"a6d430c9",
   115 => x"4966d058",
   116 => x"487129d8",
   117 => x"7098ffc3",
   118 => x"4966d07c",
   119 => x"487129d0",
   120 => x"7098ffc3",
   121 => x"4966d07c",
   122 => x"487129c8",
   123 => x"7098ffc3",
   124 => x"4866d07c",
   125 => x"7098ffc3",
   126 => x"d049757c",
   127 => x"c3487129",
   128 => x"7c7098ff",
   129 => x"f0c94b6c",
   130 => x"ffc34aff",
   131 => x"87cf05ab",
   132 => x"6c7c7149",
   133 => x"028ac14b",
   134 => x"ab7187c5",
   135 => x"7387f202",
   136 => x"264d2648",
   137 => x"264b264c",
   138 => x"49c01e4f",
   139 => x"c348d4ff",
   140 => x"81c178ff",
   141 => x"a9b7c8c3",
   142 => x"2687f104",
   143 => x"5b5e0e4f",
   144 => x"c00e5d5c",
   145 => x"f7c1f0ff",
   146 => x"c0c0c14d",
   147 => x"4bc0c0c0",
   148 => x"c487d6ff",
   149 => x"c04cdff8",
   150 => x"fd49751e",
   151 => x"86c487ce",
   152 => x"c005a8c1",
   153 => x"d4ff87e5",
   154 => x"78ffc348",
   155 => x"e1c01e73",
   156 => x"49e9c1f0",
   157 => x"c487f5fc",
   158 => x"05987086",
   159 => x"d4ff87ca",
   160 => x"78ffc348",
   161 => x"87cb48c1",
   162 => x"c187defe",
   163 => x"c6ff058c",
   164 => x"2648c087",
   165 => x"264c264d",
   166 => x"0e4f264b",
   167 => x"0e5c5b5e",
   168 => x"c1f0ffc0",
   169 => x"d4ff4cc1",
   170 => x"78ffc348",
   171 => x"f749e0cb",
   172 => x"4bd387f5",
   173 => x"49741ec0",
   174 => x"c487f1fb",
   175 => x"05987086",
   176 => x"d4ff87ca",
   177 => x"78ffc348",
   178 => x"87cb48c1",
   179 => x"c187dafd",
   180 => x"dfff058b",
   181 => x"2648c087",
   182 => x"264b264c",
   183 => x"0000004f",
   184 => x"00444d43",
   185 => x"5c5b5e0e",
   186 => x"ffc30e5d",
   187 => x"4bd4ff4d",
   188 => x"c687f6fc",
   189 => x"e1c01eea",
   190 => x"49c8c1f0",
   191 => x"c487edfa",
   192 => x"02a8c186",
   193 => x"d2fe87c8",
   194 => x"c148c087",
   195 => x"eff987e8",
   196 => x"cf497087",
   197 => x"c699ffff",
   198 => x"c802a9ea",
   199 => x"87fbfd87",
   200 => x"d1c148c0",
   201 => x"c07b7587",
   202 => x"d0fc4cf1",
   203 => x"02987087",
   204 => x"c087ecc0",
   205 => x"f0ffc01e",
   206 => x"f949fac1",
   207 => x"86c487ee",
   208 => x"da059870",
   209 => x"6b7b7587",
   210 => x"757b7549",
   211 => x"757b757b",
   212 => x"99c0c17b",
   213 => x"c187c402",
   214 => x"c087db48",
   215 => x"c287d748",
   216 => x"87ca05ac",
   217 => x"f449c0ce",
   218 => x"48c087fd",
   219 => x"8cc187c8",
   220 => x"87f6fe05",
   221 => x"4d2648c0",
   222 => x"4b264c26",
   223 => x"00004f26",
   224 => x"43484453",
   225 => x"69616620",
   226 => x"000a216c",
   227 => x"5c5b5e0e",
   228 => x"d0ff0e5d",
   229 => x"d0e5c04d",
   230 => x"c24cc0c1",
   231 => x"c148c8e1",
   232 => x"49d8d078",
   233 => x"c787c0f4",
   234 => x"f97dc24b",
   235 => x"7dc387fb",
   236 => x"49741ec0",
   237 => x"c487f5f7",
   238 => x"05a8c186",
   239 => x"c24b87c1",
   240 => x"87cb05ab",
   241 => x"f349d0d0",
   242 => x"48c087dd",
   243 => x"c187f6c0",
   244 => x"d4ff058b",
   245 => x"87ccfc87",
   246 => x"58cce1c2",
   247 => x"cd059870",
   248 => x"c01ec187",
   249 => x"d0c1f0ff",
   250 => x"87c0f749",
   251 => x"d4ff86c4",
   252 => x"78ffc348",
   253 => x"c287ccc5",
   254 => x"c258d0e1",
   255 => x"48d4ff7d",
   256 => x"c178ffc3",
   257 => x"264d2648",
   258 => x"264b264c",
   259 => x"0000004f",
   260 => x"52524549",
   261 => x"00000000",
   262 => x"00495053",
   263 => x"5c5b5e0e",
   264 => x"4d710e5d",
   265 => x"ff4cffc3",
   266 => x"7b744bd4",
   267 => x"c448d0ff",
   268 => x"7b7478c3",
   269 => x"ffc01e75",
   270 => x"49d8c1f0",
   271 => x"c487edf5",
   272 => x"02987086",
   273 => x"c8d287cb",
   274 => x"87dbf149",
   275 => x"eec048c1",
   276 => x"c37b7487",
   277 => x"c0c87bfe",
   278 => x"4966d41e",
   279 => x"c487d5f3",
   280 => x"747b7486",
   281 => x"d87b747b",
   282 => x"744ae0da",
   283 => x"c5056b7b",
   284 => x"058ac187",
   285 => x"7b7487f5",
   286 => x"c248d0ff",
   287 => x"2648c078",
   288 => x"264c264d",
   289 => x"004f264b",
   290 => x"74697257",
   291 => x"61662065",
   292 => x"64656c69",
   293 => x"5e0e000a",
   294 => x"0e5d5c5b",
   295 => x"4b7186fc",
   296 => x"c04cd4ff",
   297 => x"cdeec57e",
   298 => x"ffc34adf",
   299 => x"c3486c7c",
   300 => x"c005a8fe",
   301 => x"4d7487f8",
   302 => x"cc029b73",
   303 => x"1e66d487",
   304 => x"d2f24973",
   305 => x"d486c487",
   306 => x"48d0ff87",
   307 => x"d478d1c4",
   308 => x"ffc34a66",
   309 => x"058ac17d",
   310 => x"a6d887f8",
   311 => x"7cffc35a",
   312 => x"059b737c",
   313 => x"d0ff87c5",
   314 => x"c178d048",
   315 => x"8ac17e4a",
   316 => x"87f6fe05",
   317 => x"8efc486e",
   318 => x"4c264d26",
   319 => x"4f264b26",
   320 => x"711e731e",
   321 => x"ff4bc04a",
   322 => x"ffc348d4",
   323 => x"48d0ff78",
   324 => x"ff78c3c4",
   325 => x"ffc348d4",
   326 => x"c01e7278",
   327 => x"d1c1f0ff",
   328 => x"87c8f249",
   329 => x"987086c4",
   330 => x"c887d205",
   331 => x"66cc1ec0",
   332 => x"87e2fd49",
   333 => x"4b7086c4",
   334 => x"c248d0ff",
   335 => x"26487378",
   336 => x"0e4f264b",
   337 => x"5d5c5b5e",
   338 => x"c01ec00e",
   339 => x"c9c1f0ff",
   340 => x"87d8f149",
   341 => x"e1c21ed2",
   342 => x"f9fc49d0",
   343 => x"c086c887",
   344 => x"d284c14c",
   345 => x"f804acb7",
   346 => x"d0e1c287",
   347 => x"c349bf97",
   348 => x"c0c199c0",
   349 => x"e7c005a9",
   350 => x"d7e1c287",
   351 => x"d049bf97",
   352 => x"d8e1c231",
   353 => x"c84abf97",
   354 => x"c2b17232",
   355 => x"bf97d9e1",
   356 => x"4c71b14a",
   357 => x"ffffffcf",
   358 => x"ca84c19c",
   359 => x"87e7c134",
   360 => x"97d9e1c2",
   361 => x"31c149bf",
   362 => x"e1c299c6",
   363 => x"4abf97da",
   364 => x"722ab7c7",
   365 => x"d5e1c2b1",
   366 => x"4d4abf97",
   367 => x"e1c29dcf",
   368 => x"4abf97d6",
   369 => x"32ca9ac3",
   370 => x"97d7e1c2",
   371 => x"33c24bbf",
   372 => x"e1c2b273",
   373 => x"4bbf97d8",
   374 => x"c69bc0c3",
   375 => x"b2732bb7",
   376 => x"48c181c2",
   377 => x"49703071",
   378 => x"307548c1",
   379 => x"4c724d70",
   380 => x"947184c1",
   381 => x"adb7c0c8",
   382 => x"c187cc06",
   383 => x"c82db734",
   384 => x"01adb7c0",
   385 => x"7487f4ff",
   386 => x"264d2648",
   387 => x"264b264c",
   388 => x"5b5e0e4f",
   389 => x"f80e5d5c",
   390 => x"f8e9c286",
   391 => x"c278c048",
   392 => x"c01ef0e1",
   393 => x"87d8fb49",
   394 => x"987086c4",
   395 => x"c087c505",
   396 => x"87c0c948",
   397 => x"7ec14dc0",
   398 => x"bfdcf7c0",
   399 => x"e6e2c249",
   400 => x"4bc8714a",
   401 => x"7087dfea",
   402 => x"87c20598",
   403 => x"f7c07ec0",
   404 => x"c249bfd8",
   405 => x"714ac2e3",
   406 => x"c9ea4bc8",
   407 => x"05987087",
   408 => x"7ec087c2",
   409 => x"fdc0026e",
   410 => x"f6e8c287",
   411 => x"e9c24dbf",
   412 => x"7ebf9fee",
   413 => x"ead6c548",
   414 => x"87c705a8",
   415 => x"bff6e8c2",
   416 => x"6e87ce4d",
   417 => x"d5e9ca48",
   418 => x"87c502a8",
   419 => x"e3c748c0",
   420 => x"f0e1c287",
   421 => x"f949751e",
   422 => x"86c487e6",
   423 => x"c5059870",
   424 => x"c748c087",
   425 => x"f7c087ce",
   426 => x"c249bfd8",
   427 => x"714ac2e3",
   428 => x"f1e84bc8",
   429 => x"05987087",
   430 => x"e9c287c8",
   431 => x"78c148f8",
   432 => x"f7c087da",
   433 => x"c249bfdc",
   434 => x"714ae6e2",
   435 => x"d5e84bc8",
   436 => x"02987087",
   437 => x"c087c5c0",
   438 => x"87d8c648",
   439 => x"97eee9c2",
   440 => x"d5c149bf",
   441 => x"cdc005a9",
   442 => x"efe9c287",
   443 => x"c249bf97",
   444 => x"c002a9ea",
   445 => x"48c087c5",
   446 => x"c287f9c5",
   447 => x"bf97f0e1",
   448 => x"e9c3487e",
   449 => x"cec002a8",
   450 => x"c3486e87",
   451 => x"c002a8eb",
   452 => x"48c087c5",
   453 => x"c287ddc5",
   454 => x"bf97fbe1",
   455 => x"c0059949",
   456 => x"e1c287cc",
   457 => x"49bf97fc",
   458 => x"c002a9c2",
   459 => x"48c087c5",
   460 => x"c287c1c5",
   461 => x"bf97fde1",
   462 => x"f4e9c248",
   463 => x"484c7058",
   464 => x"e9c288c1",
   465 => x"e1c258f8",
   466 => x"49bf97fe",
   467 => x"e1c28175",
   468 => x"4abf97ff",
   469 => x"a17232c8",
   470 => x"c8eec27e",
   471 => x"c2786e48",
   472 => x"bf97c0e2",
   473 => x"58a6c848",
   474 => x"bff8e9c2",
   475 => x"87cfc202",
   476 => x"bfd8f7c0",
   477 => x"c2e3c249",
   478 => x"4bc8714a",
   479 => x"7087e7e5",
   480 => x"c5c00298",
   481 => x"c348c087",
   482 => x"e9c287ea",
   483 => x"c24cbff0",
   484 => x"c25cdcee",
   485 => x"bf97d5e2",
   486 => x"c231c849",
   487 => x"bf97d4e2",
   488 => x"c249a14a",
   489 => x"bf97d6e2",
   490 => x"7232d04a",
   491 => x"e2c249a1",
   492 => x"4abf97d7",
   493 => x"a17232d8",
   494 => x"9166c449",
   495 => x"bfc8eec2",
   496 => x"d0eec281",
   497 => x"dde2c259",
   498 => x"c84abf97",
   499 => x"dce2c232",
   500 => x"a24bbf97",
   501 => x"dee2c24a",
   502 => x"d04bbf97",
   503 => x"4aa27333",
   504 => x"97dfe2c2",
   505 => x"9bcf4bbf",
   506 => x"a27333d8",
   507 => x"d4eec24a",
   508 => x"748ac25a",
   509 => x"d4eec292",
   510 => x"78a17248",
   511 => x"c287c1c1",
   512 => x"bf97c2e2",
   513 => x"c231c849",
   514 => x"bf97c1e2",
   515 => x"c549a14a",
   516 => x"81ffc731",
   517 => x"eec229c9",
   518 => x"e2c259dc",
   519 => x"4abf97c7",
   520 => x"e2c232c8",
   521 => x"4bbf97c6",
   522 => x"66c44aa2",
   523 => x"c2826e92",
   524 => x"c25ad8ee",
   525 => x"c048d0ee",
   526 => x"cceec278",
   527 => x"78a17248",
   528 => x"48dceec2",
   529 => x"bfd0eec2",
   530 => x"e0eec278",
   531 => x"d4eec248",
   532 => x"e9c278bf",
   533 => x"c002bff8",
   534 => x"487487c9",
   535 => x"7e7030c4",
   536 => x"c287c9c0",
   537 => x"48bfd8ee",
   538 => x"7e7030c4",
   539 => x"48fce9c2",
   540 => x"48c1786e",
   541 => x"4d268ef8",
   542 => x"4b264c26",
   543 => x"5e0e4f26",
   544 => x"0e5d5c5b",
   545 => x"e9c24a71",
   546 => x"cb02bff8",
   547 => x"c74b7287",
   548 => x"c14d722b",
   549 => x"87c99dff",
   550 => x"2bc84b72",
   551 => x"ffc34d72",
   552 => x"c8eec29d",
   553 => x"f7c083bf",
   554 => x"02abbfd4",
   555 => x"f7c087d9",
   556 => x"e1c25bd8",
   557 => x"49731ef0",
   558 => x"c487c5f1",
   559 => x"05987086",
   560 => x"48c087c5",
   561 => x"c287e6c0",
   562 => x"02bff8e9",
   563 => x"497587d2",
   564 => x"e1c291c4",
   565 => x"4c6981f0",
   566 => x"ffffffcf",
   567 => x"87cb9cff",
   568 => x"91c24975",
   569 => x"81f0e1c2",
   570 => x"744c699f",
   571 => x"264d2648",
   572 => x"264b264c",
   573 => x"5b5e0e4f",
   574 => x"f40e5d5c",
   575 => x"59a6cc86",
   576 => x"c50566c8",
   577 => x"c348c087",
   578 => x"66c887c8",
   579 => x"7080c848",
   580 => x"78c0487e",
   581 => x"c70266dc",
   582 => x"9766dc87",
   583 => x"87c505bf",
   584 => x"edc248c0",
   585 => x"c11ec087",
   586 => x"eeca4949",
   587 => x"7086c487",
   588 => x"c0029c4c",
   589 => x"eac287fc",
   590 => x"66dc4ac0",
   591 => x"cadeff49",
   592 => x"02987087",
   593 => x"7487ebc0",
   594 => x"4966dc4a",
   595 => x"deff4bcb",
   596 => x"987087ee",
   597 => x"c087db02",
   598 => x"029c741e",
   599 => x"4dc087c4",
   600 => x"4dc187c2",
   601 => x"f2c94975",
   602 => x"7086c487",
   603 => x"ff059c4c",
   604 => x"9c7487c4",
   605 => x"87d8c102",
   606 => x"6e49a4dc",
   607 => x"da786948",
   608 => x"66c849a4",
   609 => x"c880c448",
   610 => x"699f58a6",
   611 => x"0866c448",
   612 => x"f8e9c278",
   613 => x"87d202bf",
   614 => x"9f49a4d4",
   615 => x"ffc04969",
   616 => x"487199ff",
   617 => x"7e7030d0",
   618 => x"7ec087c2",
   619 => x"c448496e",
   620 => x"c480bf66",
   621 => x"c8780866",
   622 => x"78c04866",
   623 => x"cc4966c8",
   624 => x"bf66c481",
   625 => x"4966c879",
   626 => x"79c081d0",
   627 => x"87c248c1",
   628 => x"8ef448c0",
   629 => x"4c264d26",
   630 => x"4f264b26",
   631 => x"5c5b5e0e",
   632 => x"4c710e5d",
   633 => x"744d66d0",
   634 => x"c6c1029c",
   635 => x"49a4c887",
   636 => x"fec00269",
   637 => x"6c4a7587",
   638 => x"4da17249",
   639 => x"f4e9c2b9",
   640 => x"baff4abf",
   641 => x"99719972",
   642 => x"87e5c002",
   643 => x"6b4ba4c4",
   644 => x"87eaf949",
   645 => x"e9c27b70",
   646 => x"6c49bff0",
   647 => x"757c7181",
   648 => x"e9c2b94a",
   649 => x"ff4abff4",
   650 => x"719972ba",
   651 => x"dbff0599",
   652 => x"267c7587",
   653 => x"264c264d",
   654 => x"1e4f264b",
   655 => x"4b711e73",
   656 => x"87c7029b",
   657 => x"6949a3c8",
   658 => x"c087c505",
   659 => x"87f6c048",
   660 => x"bfcceec2",
   661 => x"4aa3c449",
   662 => x"8ac24a6a",
   663 => x"bff0e9c2",
   664 => x"49a17292",
   665 => x"bff4e9c2",
   666 => x"729a6b4a",
   667 => x"f7c049a1",
   668 => x"66c859d8",
   669 => x"c7ea711e",
   670 => x"7086c487",
   671 => x"87c40598",
   672 => x"87c248c0",
   673 => x"4b2648c1",
   674 => x"731e4f26",
   675 => x"9b4b711e",
   676 => x"c887c702",
   677 => x"056949a3",
   678 => x"48c087c5",
   679 => x"c287f6c0",
   680 => x"49bfccee",
   681 => x"6a4aa3c4",
   682 => x"c28ac24a",
   683 => x"92bff0e9",
   684 => x"c249a172",
   685 => x"4abff4e9",
   686 => x"a1729a6b",
   687 => x"d8f7c049",
   688 => x"1e66c859",
   689 => x"87d4e571",
   690 => x"987086c4",
   691 => x"c087c405",
   692 => x"c187c248",
   693 => x"264b2648",
   694 => x"5b5e0e4f",
   695 => x"fc0e5d5c",
   696 => x"d44b7186",
   697 => x"9b734d66",
   698 => x"87ccc102",
   699 => x"6949a3c8",
   700 => x"87c4c102",
   701 => x"c24ca3d0",
   702 => x"49bff4e9",
   703 => x"4a6cb9ff",
   704 => x"66d47e99",
   705 => x"87cd06a9",
   706 => x"cc7c7bc0",
   707 => x"a3c44aa3",
   708 => x"ca796a49",
   709 => x"f8497287",
   710 => x"66d499c0",
   711 => x"758d714d",
   712 => x"7129c949",
   713 => x"fa49731e",
   714 => x"e1c287f2",
   715 => x"49731ef0",
   716 => x"c887c8fc",
   717 => x"7c66d486",
   718 => x"4d268efc",
   719 => x"4b264c26",
   720 => x"731e4f26",
   721 => x"9b4b711e",
   722 => x"87e4c002",
   723 => x"5be0eec2",
   724 => x"8ac24a73",
   725 => x"bff0e9c2",
   726 => x"eec29249",
   727 => x"7248bfcc",
   728 => x"e4eec280",
   729 => x"c4487158",
   730 => x"c0eac230",
   731 => x"87edc058",
   732 => x"48dceec2",
   733 => x"bfd0eec2",
   734 => x"e0eec278",
   735 => x"d4eec248",
   736 => x"e9c278bf",
   737 => x"c902bff8",
   738 => x"f0e9c287",
   739 => x"31c449bf",
   740 => x"eec287c7",
   741 => x"c449bfd8",
   742 => x"c0eac231",
   743 => x"264b2659",
   744 => x"5b5e0e4f",
   745 => x"4a710e5c",
   746 => x"9a724bc0",
   747 => x"87e0c002",
   748 => x"9f49a2da",
   749 => x"e9c24b69",
   750 => x"cf02bff8",
   751 => x"49a2d487",
   752 => x"4c49699f",
   753 => x"9cffffc0",
   754 => x"87c234d0",
   755 => x"b3744cc0",
   756 => x"edfd4973",
   757 => x"264c2687",
   758 => x"0e4f264b",
   759 => x"5d5c5b5e",
   760 => x"c886f00e",
   761 => x"ffcf59a6",
   762 => x"4cf8ffff",
   763 => x"66c47ec0",
   764 => x"c287d802",
   765 => x"c048ece1",
   766 => x"e4e1c278",
   767 => x"e0eec248",
   768 => x"e1c278bf",
   769 => x"eec248e8",
   770 => x"c278bfdc",
   771 => x"c048cdea",
   772 => x"fce9c250",
   773 => x"e1c249bf",
   774 => x"714abfec",
   775 => x"cbc403aa",
   776 => x"cf497287",
   777 => x"e9c00599",
   778 => x"d4f7c087",
   779 => x"e4e1c248",
   780 => x"e1c278bf",
   781 => x"e1c21ef0",
   782 => x"c249bfe4",
   783 => x"c148e4e1",
   784 => x"e27178a1",
   785 => x"86c487fa",
   786 => x"48d0f7c0",
   787 => x"78f0e1c2",
   788 => x"f7c087cc",
   789 => x"c048bfd0",
   790 => x"f7c080e0",
   791 => x"e1c258d4",
   792 => x"c148bfec",
   793 => x"f0e1c280",
   794 => x"0dd02758",
   795 => x"97bf0000",
   796 => x"029d4dbf",
   797 => x"c387e5c2",
   798 => x"c202ade5",
   799 => x"f7c087de",
   800 => x"cb4bbfd0",
   801 => x"4c1149a3",
   802 => x"c105accf",
   803 => x"497587d2",
   804 => x"89c199df",
   805 => x"eac291cd",
   806 => x"a3c181c0",
   807 => x"c351124a",
   808 => x"51124aa3",
   809 => x"124aa3c5",
   810 => x"4aa3c751",
   811 => x"a3c95112",
   812 => x"ce51124a",
   813 => x"51124aa3",
   814 => x"124aa3d0",
   815 => x"4aa3d251",
   816 => x"a3d45112",
   817 => x"d651124a",
   818 => x"51124aa3",
   819 => x"124aa3d8",
   820 => x"4aa3dc51",
   821 => x"a3de5112",
   822 => x"c151124a",
   823 => x"87fcc07e",
   824 => x"99c84974",
   825 => x"87edc005",
   826 => x"99d04974",
   827 => x"c087d305",
   828 => x"c00266e0",
   829 => x"497387cc",
   830 => x"0f66e0c0",
   831 => x"c0029870",
   832 => x"056e87d3",
   833 => x"c287c6c0",
   834 => x"c048c0ea",
   835 => x"d0f7c050",
   836 => x"ebc248bf",
   837 => x"cdeac287",
   838 => x"7e50c048",
   839 => x"bffce9c2",
   840 => x"ece1c249",
   841 => x"aa714abf",
   842 => x"87f5fb04",
   843 => x"ffffffcf",
   844 => x"eec24cf8",
   845 => x"c005bfe0",
   846 => x"e9c287c8",
   847 => x"c102bff8",
   848 => x"e1c287fc",
   849 => x"ec49bfe8",
   850 => x"e1c287f4",
   851 => x"a6c458ec",
   852 => x"e8e1c248",
   853 => x"e9c278bf",
   854 => x"c002bff8",
   855 => x"66c487db",
   856 => x"74997449",
   857 => x"c8c002a9",
   858 => x"48a6c887",
   859 => x"e7c078c0",
   860 => x"48a6c887",
   861 => x"dfc078c1",
   862 => x"4966c487",
   863 => x"99f8ffcf",
   864 => x"c8c002a9",
   865 => x"48a6cc87",
   866 => x"c5c078c0",
   867 => x"48a6cc87",
   868 => x"a6c878c1",
   869 => x"7866cc48",
   870 => x"c00566c8",
   871 => x"66c487e0",
   872 => x"c289c249",
   873 => x"4abff0e9",
   874 => x"cceec291",
   875 => x"e1c24abf",
   876 => x"a17248e4",
   877 => x"ece1c278",
   878 => x"f978c048",
   879 => x"48c087d3",
   880 => x"ffffffcf",
   881 => x"8ef04cf8",
   882 => x"4c264d26",
   883 => x"4f264b26",
   884 => x"00000000",
   885 => x"ffffffff",
   886 => x"00000de0",
   887 => x"00000dec",
   888 => x"33544146",
   889 => x"20202032",
   890 => x"00000000",
   891 => x"31544146",
   892 => x"20202036",
   893 => x"d4ff1e00",
   894 => x"78ffc348",
   895 => x"4f264868",
   896 => x"48d4ff1e",
   897 => x"ff78ffc3",
   898 => x"e1c048d0",
   899 => x"48d4ff78",
   900 => x"4f2678d4",
   901 => x"48d0ff1e",
   902 => x"2678e0c0",
   903 => x"d4ff1e4f",
   904 => x"99497087",
   905 => x"c087c602",
   906 => x"f105a9fb",
   907 => x"26487187",
   908 => x"5b5e0e4f",
   909 => x"4b710e5c",
   910 => x"f8fe4cc0",
   911 => x"99497087",
   912 => x"87f9c002",
   913 => x"02a9ecc0",
   914 => x"c087f2c0",
   915 => x"c002a9fb",
   916 => x"66cc87eb",
   917 => x"c703acb7",
   918 => x"0266d087",
   919 => x"537187c2",
   920 => x"c2029971",
   921 => x"fe84c187",
   922 => x"497087cb",
   923 => x"87cd0299",
   924 => x"02a9ecc0",
   925 => x"fbc087c7",
   926 => x"d5ff05a9",
   927 => x"0266d087",
   928 => x"97c087c3",
   929 => x"a9ecc07b",
   930 => x"7487c405",
   931 => x"7487c54a",
   932 => x"8a0ac04a",
   933 => x"4c264872",
   934 => x"4f264b26",
   935 => x"87d5fd1e",
   936 => x"c04a4970",
   937 => x"c904aaf0",
   938 => x"aaf9c087",
   939 => x"c087c301",
   940 => x"c1c18af0",
   941 => x"87c904aa",
   942 => x"01aadac1",
   943 => x"f7c087c3",
   944 => x"2648728a",
   945 => x"5b5e0e4f",
   946 => x"f80e5d5c",
   947 => x"c04c7186",
   948 => x"87ecfc7e",
   949 => x"fdc04bc0",
   950 => x"49bf97e4",
   951 => x"cf04a9c0",
   952 => x"87f9fc87",
   953 => x"fdc083c1",
   954 => x"49bf97e4",
   955 => x"87f106ab",
   956 => x"97e4fdc0",
   957 => x"87cf02bf",
   958 => x"7087fafb",
   959 => x"c6029949",
   960 => x"a9ecc087",
   961 => x"c087f105",
   962 => x"87e9fb4b",
   963 => x"e4fb4d70",
   964 => x"58a6c887",
   965 => x"7087defb",
   966 => x"c883c14a",
   967 => x"699749a4",
   968 => x"da05ad49",
   969 => x"49a4c987",
   970 => x"c4496997",
   971 => x"ce05a966",
   972 => x"49a4ca87",
   973 => x"aa496997",
   974 => x"c187c405",
   975 => x"c087d07e",
   976 => x"c602adec",
   977 => x"adfbc087",
   978 => x"c087c405",
   979 => x"6e7ec14b",
   980 => x"87f5fe02",
   981 => x"7387fdfa",
   982 => x"268ef848",
   983 => x"264c264d",
   984 => x"004f264b",
   985 => x"1e731e00",
   986 => x"c84bd4ff",
   987 => x"d0ff4a66",
   988 => x"78c5c848",
   989 => x"c148d4ff",
   990 => x"7b1178d4",
   991 => x"f9058ac1",
   992 => x"48d0ff87",
   993 => x"4b2678c4",
   994 => x"5e0e4f26",
   995 => x"0e5d5c5b",
   996 => x"7e7186f8",
   997 => x"eec21e6e",
   998 => x"d8e549f0",
   999 => x"7086c487",
  1000 => x"e4c40298",
  1001 => x"e0edc187",
  1002 => x"496e4cbf",
  1003 => x"c887d6fc",
  1004 => x"987058a6",
  1005 => x"c487c505",
  1006 => x"78c148a6",
  1007 => x"c548d0ff",
  1008 => x"48d4ff78",
  1009 => x"c478d5c1",
  1010 => x"89c14966",
  1011 => x"edc131c6",
  1012 => x"4abf97d8",
  1013 => x"ffb07148",
  1014 => x"ff7808d4",
  1015 => x"78c448d0",
  1016 => x"97eceec2",
  1017 => x"99d049bf",
  1018 => x"c587dd02",
  1019 => x"48d4ff78",
  1020 => x"c078d6c1",
  1021 => x"48d4ff4a",
  1022 => x"c178ffc3",
  1023 => x"aae0c082",
  1024 => x"ff87f204",
  1025 => x"78c448d0",
  1026 => x"c348d4ff",
  1027 => x"d0ff78ff",
  1028 => x"ff78c548",
  1029 => x"d3c148d4",
  1030 => x"ff78c178",
  1031 => x"78c448d0",
  1032 => x"06acb7c0",
  1033 => x"c287cbc2",
  1034 => x"4bbff8ee",
  1035 => x"737e748c",
  1036 => x"ddc1029b",
  1037 => x"4dc0c887",
  1038 => x"abb7c08b",
  1039 => x"c887c603",
  1040 => x"c04da3c0",
  1041 => x"eceec24b",
  1042 => x"d049bf97",
  1043 => x"87cf0299",
  1044 => x"eec21ec0",
  1045 => x"e2e749f0",
  1046 => x"7086c487",
  1047 => x"c287d84c",
  1048 => x"c21ef0e1",
  1049 => x"e749f0ee",
  1050 => x"4c7087d1",
  1051 => x"e1c21e75",
  1052 => x"f0fb49f0",
  1053 => x"7486c887",
  1054 => x"87c5059c",
  1055 => x"cac148c0",
  1056 => x"c21ec187",
  1057 => x"e549f0ee",
  1058 => x"86c487d2",
  1059 => x"fe059b73",
  1060 => x"4c6e87e3",
  1061 => x"06acb7c0",
  1062 => x"eec287d1",
  1063 => x"78c048f0",
  1064 => x"78c080d0",
  1065 => x"eec280f4",
  1066 => x"c078bffc",
  1067 => x"fd01acb7",
  1068 => x"d0ff87f5",
  1069 => x"ff78c548",
  1070 => x"d3c148d4",
  1071 => x"ff78c078",
  1072 => x"78c448d0",
  1073 => x"c2c048c1",
  1074 => x"f848c087",
  1075 => x"264d268e",
  1076 => x"264b264c",
  1077 => x"5b5e0e4f",
  1078 => x"fc0e5d5c",
  1079 => x"c04d7186",
  1080 => x"04ad4c4b",
  1081 => x"c087e8c0",
  1082 => x"741ec5fb",
  1083 => x"87c4029c",
  1084 => x"87c24ac0",
  1085 => x"49724ac1",
  1086 => x"c487e0eb",
  1087 => x"c17e7086",
  1088 => x"c2056e83",
  1089 => x"c14b7587",
  1090 => x"06ab7584",
  1091 => x"6e87d8ff",
  1092 => x"268efc48",
  1093 => x"264c264d",
  1094 => x"0e4f264b",
  1095 => x"0e5c5b5e",
  1096 => x"66cc4b71",
  1097 => x"4c87d802",
  1098 => x"028cf0c0",
  1099 => x"4a7487d8",
  1100 => x"d1028ac1",
  1101 => x"cd028a87",
  1102 => x"c9028a87",
  1103 => x"7387d987",
  1104 => x"87c6f949",
  1105 => x"1e7487d2",
  1106 => x"d9c149c0",
  1107 => x"1e7487f2",
  1108 => x"d9c14973",
  1109 => x"86c887ea",
  1110 => x"4b264c26",
  1111 => x"5e0e4f26",
  1112 => x"0e5d5c5b",
  1113 => x"4c7186fc",
  1114 => x"c291de49",
  1115 => x"714ddcef",
  1116 => x"026d9785",
  1117 => x"c287dcc1",
  1118 => x"49bfccef",
  1119 => x"fd718174",
  1120 => x"7e7087d3",
  1121 => x"c0029848",
  1122 => x"efc287f2",
  1123 => x"4a704bd0",
  1124 => x"fefe49cb",
  1125 => x"4b7487ce",
  1126 => x"edc193cc",
  1127 => x"83c483e4",
  1128 => x"7be0c7c1",
  1129 => x"c4c14974",
  1130 => x"7b7587e2",
  1131 => x"97dcedc1",
  1132 => x"c21e49bf",
  1133 => x"fd49d0ef",
  1134 => x"86c487e1",
  1135 => x"c4c14974",
  1136 => x"49c087ca",
  1137 => x"87e5c5c1",
  1138 => x"48e8eec2",
  1139 => x"c04950c0",
  1140 => x"fc87cce2",
  1141 => x"264d268e",
  1142 => x"264b264c",
  1143 => x"0000004f",
  1144 => x"64616f4c",
  1145 => x"2e676e69",
  1146 => x"1e002e2e",
  1147 => x"4b711e73",
  1148 => x"ccefc249",
  1149 => x"fb7181bf",
  1150 => x"4a7087db",
  1151 => x"87c4029a",
  1152 => x"87dde649",
  1153 => x"48ccefc2",
  1154 => x"497378c0",
  1155 => x"2687fac1",
  1156 => x"1e4f264b",
  1157 => x"4b711e73",
  1158 => x"024aa3c4",
  1159 => x"c187d0c1",
  1160 => x"87dc028a",
  1161 => x"f2c0028a",
  1162 => x"c1058a87",
  1163 => x"efc287d3",
  1164 => x"c102bfcc",
  1165 => x"c14887cb",
  1166 => x"d0efc288",
  1167 => x"87c1c158",
  1168 => x"bfccefc2",
  1169 => x"c289c649",
  1170 => x"c059d0ef",
  1171 => x"c003a9b7",
  1172 => x"efc287ef",
  1173 => x"78c048cc",
  1174 => x"c287e6c0",
  1175 => x"02bfc8ef",
  1176 => x"efc287df",
  1177 => x"c148bfcc",
  1178 => x"d0efc280",
  1179 => x"c287d258",
  1180 => x"02bfc8ef",
  1181 => x"efc287cb",
  1182 => x"c648bfcc",
  1183 => x"d0efc280",
  1184 => x"c4497358",
  1185 => x"264b2687",
  1186 => x"5b5e0e4f",
  1187 => x"f00e5d5c",
  1188 => x"59a6d086",
  1189 => x"4df0e1c2",
  1190 => x"efc24cc0",
  1191 => x"78c148c8",
  1192 => x"c048a6c4",
  1193 => x"c27e7578",
  1194 => x"48bfccef",
  1195 => x"c006a8c0",
  1196 => x"7e7587fa",
  1197 => x"48f0e1c2",
  1198 => x"efc00298",
  1199 => x"c5fbc087",
  1200 => x"0266c81e",
  1201 => x"4dc087c4",
  1202 => x"4dc187c2",
  1203 => x"cae44975",
  1204 => x"7086c487",
  1205 => x"c484c17e",
  1206 => x"80c14866",
  1207 => x"c258a6c8",
  1208 => x"acbfccef",
  1209 => x"6e87c503",
  1210 => x"87d1ff05",
  1211 => x"4cc04d6e",
  1212 => x"c3029d75",
  1213 => x"fbc087e0",
  1214 => x"66c81ec5",
  1215 => x"cc87c702",
  1216 => x"78c048a6",
  1217 => x"a6cc87c5",
  1218 => x"cc78c148",
  1219 => x"cae34966",
  1220 => x"7086c487",
  1221 => x"0298487e",
  1222 => x"4987e8c2",
  1223 => x"699781cb",
  1224 => x"0299d049",
  1225 => x"c187d6c1",
  1226 => x"744aebc7",
  1227 => x"c191cc49",
  1228 => x"7281e4ed",
  1229 => x"c381c879",
  1230 => x"497451ff",
  1231 => x"efc291de",
  1232 => x"85714ddc",
  1233 => x"7d97c1c2",
  1234 => x"c049a5c1",
  1235 => x"eac251e0",
  1236 => x"02bf97c0",
  1237 => x"84c187d2",
  1238 => x"c24ba5c2",
  1239 => x"db4ac0ea",
  1240 => x"fff6fe49",
  1241 => x"87dbc187",
  1242 => x"c049a5cd",
  1243 => x"c284c151",
  1244 => x"4a6e4ba5",
  1245 => x"f6fe49cb",
  1246 => x"c6c187ea",
  1247 => x"dec5c187",
  1248 => x"cc49744a",
  1249 => x"e4edc191",
  1250 => x"c2797281",
  1251 => x"bf97c0ea",
  1252 => x"7487d802",
  1253 => x"c191de49",
  1254 => x"dcefc284",
  1255 => x"c283714b",
  1256 => x"dd4ac0ea",
  1257 => x"fbf5fe49",
  1258 => x"7487d887",
  1259 => x"c293de4b",
  1260 => x"cb83dcef",
  1261 => x"51c049a3",
  1262 => x"6e7384c1",
  1263 => x"fe49cb4a",
  1264 => x"c487e1f5",
  1265 => x"80c14866",
  1266 => x"c758a6c8",
  1267 => x"c5c003ac",
  1268 => x"fc056e87",
  1269 => x"acc787e0",
  1270 => x"87e6c003",
  1271 => x"48c8efc2",
  1272 => x"c5c178c0",
  1273 => x"49744ade",
  1274 => x"edc191cc",
  1275 => x"797281e4",
  1276 => x"91de4974",
  1277 => x"81dcefc2",
  1278 => x"84c151c0",
  1279 => x"ff04acc7",
  1280 => x"efc187da",
  1281 => x"50c048c0",
  1282 => x"d1c180f7",
  1283 => x"d0c140f9",
  1284 => x"80c878ec",
  1285 => x"78d3c8c1",
  1286 => x"c04966cc",
  1287 => x"f087edfa",
  1288 => x"264d268e",
  1289 => x"264b264c",
  1290 => x"0000004f",
  1291 => x"61422080",
  1292 => x"1e006b63",
  1293 => x"4b711e73",
  1294 => x"c191cc49",
  1295 => x"c881e4ed",
  1296 => x"edc14aa1",
  1297 => x"501248d8",
  1298 => x"c04aa1c9",
  1299 => x"1248e4fd",
  1300 => x"c181ca50",
  1301 => x"1148dced",
  1302 => x"dcedc150",
  1303 => x"1e49bf97",
  1304 => x"f6f249c0",
  1305 => x"f8497387",
  1306 => x"8efc87df",
  1307 => x"4f264b26",
  1308 => x"c049c01e",
  1309 => x"2687f6fa",
  1310 => x"4a711e4f",
  1311 => x"c191cc49",
  1312 => x"c881e4ed",
  1313 => x"e8eec281",
  1314 => x"c0501148",
  1315 => x"fe49a2f0",
  1316 => x"c087f9ef",
  1317 => x"87c7d749",
  1318 => x"ff1e4f26",
  1319 => x"ffc34ad4",
  1320 => x"48d0ff7a",
  1321 => x"de78e1c0",
  1322 => x"487a717a",
  1323 => x"7028b7c8",
  1324 => x"d048717a",
  1325 => x"7a7028b7",
  1326 => x"b7d84871",
  1327 => x"ff7a7028",
  1328 => x"e0c048d0",
  1329 => x"0e4f2678",
  1330 => x"5d5c5b5e",
  1331 => x"7186f40e",
  1332 => x"91cc494d",
  1333 => x"81e4edc1",
  1334 => x"ca4aa1c8",
  1335 => x"a6c47ea1",
  1336 => x"e4eec248",
  1337 => x"976e78bf",
  1338 => x"66c44bbf",
  1339 => x"122c734c",
  1340 => x"58a6cc48",
  1341 => x"84c19c70",
  1342 => x"699781c9",
  1343 => x"04acb749",
  1344 => x"4cc087c2",
  1345 => x"4abf976e",
  1346 => x"724966c8",
  1347 => x"c4b9ff31",
  1348 => x"48749966",
  1349 => x"4a703072",
  1350 => x"e8eec2b1",
  1351 => x"f9fd7159",
  1352 => x"c21ec787",
  1353 => x"1ebfc4ef",
  1354 => x"1ee4edc1",
  1355 => x"97e8eec2",
  1356 => x"f4c149bf",
  1357 => x"c0497587",
  1358 => x"e887d1f6",
  1359 => x"264d268e",
  1360 => x"264b264c",
  1361 => x"1e731e4f",
  1362 => x"fd494b71",
  1363 => x"497387f9",
  1364 => x"2687f4fd",
  1365 => x"1e4f264b",
  1366 => x"4b711e73",
  1367 => x"024aa3c2",
  1368 => x"8ac187d6",
  1369 => x"87e2c005",
  1370 => x"bfc4efc2",
  1371 => x"4887db02",
  1372 => x"efc288c1",
  1373 => x"87d258c8",
  1374 => x"bfc8efc2",
  1375 => x"c287cb02",
  1376 => x"48bfc4ef",
  1377 => x"efc280c1",
  1378 => x"1ec758c8",
  1379 => x"bfc4efc2",
  1380 => x"e4edc11e",
  1381 => x"e8eec21e",
  1382 => x"cc49bf97",
  1383 => x"c0497387",
  1384 => x"f487e9f4",
  1385 => x"264b268e",
  1386 => x"5b5e0e4f",
  1387 => x"ff0e5d5c",
  1388 => x"e4c086cc",
  1389 => x"a6cc59a6",
  1390 => x"c478c048",
  1391 => x"c478c080",
  1392 => x"66c8c180",
  1393 => x"c180c478",
  1394 => x"c180c478",
  1395 => x"c8efc278",
  1396 => x"e078c148",
  1397 => x"c4e187ea",
  1398 => x"87d9e087",
  1399 => x"fbc04c70",
  1400 => x"f3c102ac",
  1401 => x"66e0c087",
  1402 => x"87e8c105",
  1403 => x"4a66c4c1",
  1404 => x"7e6a82c4",
  1405 => x"48c0e9c1",
  1406 => x"4120496e",
  1407 => x"51104120",
  1408 => x"4866c4c1",
  1409 => x"78f3d0c1",
  1410 => x"81c7496a",
  1411 => x"c4c15174",
  1412 => x"81c84966",
  1413 => x"a6d851c1",
  1414 => x"c178c248",
  1415 => x"c94966c4",
  1416 => x"c151c081",
  1417 => x"ca4966c4",
  1418 => x"c151c081",
  1419 => x"6a1ed81e",
  1420 => x"ff81c849",
  1421 => x"c887fadf",
  1422 => x"66c8c186",
  1423 => x"01a8c048",
  1424 => x"a6d087c7",
  1425 => x"cf78c148",
  1426 => x"66c8c187",
  1427 => x"d888c148",
  1428 => x"87c458a6",
  1429 => x"87c5dfff",
  1430 => x"cd029c74",
  1431 => x"66d087da",
  1432 => x"66ccc148",
  1433 => x"cfcd03a8",
  1434 => x"48a6c887",
  1435 => x"ff7e78c0",
  1436 => x"7087c2de",
  1437 => x"acd0c14c",
  1438 => x"87e7c205",
  1439 => x"6e48a6c4",
  1440 => x"87d8e078",
  1441 => x"cc487e70",
  1442 => x"c506a866",
  1443 => x"48a6cc87",
  1444 => x"ddff786e",
  1445 => x"4c7087df",
  1446 => x"05acecc0",
  1447 => x"d087eec1",
  1448 => x"91cc4966",
  1449 => x"8166c4c1",
  1450 => x"6a4aa1c4",
  1451 => x"4aa1c84d",
  1452 => x"d1c1526e",
  1453 => x"dcff79f9",
  1454 => x"4c7087fb",
  1455 => x"87d9029c",
  1456 => x"02acfbc0",
  1457 => x"557487d3",
  1458 => x"87e9dcff",
  1459 => x"029c4c70",
  1460 => x"fbc087c7",
  1461 => x"edff05ac",
  1462 => x"55e0c087",
  1463 => x"c055c1c2",
  1464 => x"e0c07d97",
  1465 => x"66c44866",
  1466 => x"87db05a8",
  1467 => x"d44866d0",
  1468 => x"ca04a866",
  1469 => x"4866d087",
  1470 => x"a6d480c1",
  1471 => x"d487c858",
  1472 => x"88c14866",
  1473 => x"ff58a6d8",
  1474 => x"7087eadb",
  1475 => x"acd0c14c",
  1476 => x"dc87c905",
  1477 => x"80c14866",
  1478 => x"58a6e0c0",
  1479 => x"02acd0c1",
  1480 => x"6e87d9fd",
  1481 => x"66e0c048",
  1482 => x"ebc905a8",
  1483 => x"a6e4c087",
  1484 => x"7478c048",
  1485 => x"88fbc048",
  1486 => x"7058a6c8",
  1487 => x"ddc90298",
  1488 => x"88cb4887",
  1489 => x"7058a6c8",
  1490 => x"cfc10298",
  1491 => x"88c94887",
  1492 => x"7058a6c8",
  1493 => x"ffc30298",
  1494 => x"88c44887",
  1495 => x"7058a6c8",
  1496 => x"87cf0298",
  1497 => x"c888c148",
  1498 => x"987058a6",
  1499 => x"87e8c302",
  1500 => x"c887dcc8",
  1501 => x"f0c048a6",
  1502 => x"f8d9ff78",
  1503 => x"c04c7087",
  1504 => x"c002acec",
  1505 => x"a6cc87c3",
  1506 => x"acecc05c",
  1507 => x"ff87cd02",
  1508 => x"7087e2d9",
  1509 => x"acecc04c",
  1510 => x"87f3ff05",
  1511 => x"02acecc0",
  1512 => x"ff87c4c0",
  1513 => x"c087ced9",
  1514 => x"d81eca1e",
  1515 => x"91cc4966",
  1516 => x"4866ccc1",
  1517 => x"a6cc8071",
  1518 => x"4866c858",
  1519 => x"a6d080c4",
  1520 => x"bf66cc58",
  1521 => x"e8d9ff49",
  1522 => x"de1ec187",
  1523 => x"bf66d41e",
  1524 => x"dcd9ff49",
  1525 => x"7086d087",
  1526 => x"08c04849",
  1527 => x"a6ecc088",
  1528 => x"06a8c058",
  1529 => x"c087eec0",
  1530 => x"dd4866e8",
  1531 => x"e4c003a8",
  1532 => x"bf66c487",
  1533 => x"66e8c049",
  1534 => x"51e0c081",
  1535 => x"4966e8c0",
  1536 => x"66c481c1",
  1537 => x"c1c281bf",
  1538 => x"66e8c051",
  1539 => x"c481c249",
  1540 => x"c081bf66",
  1541 => x"c1486e51",
  1542 => x"6e78f3d0",
  1543 => x"d881c849",
  1544 => x"496e5166",
  1545 => x"66dc81c9",
  1546 => x"ca496e51",
  1547 => x"5166c881",
  1548 => x"c14866d8",
  1549 => x"58a6dc80",
  1550 => x"d44866d0",
  1551 => x"c004a866",
  1552 => x"66d087cb",
  1553 => x"d480c148",
  1554 => x"d1c558a6",
  1555 => x"4866d487",
  1556 => x"a6d888c1",
  1557 => x"87c6c558",
  1558 => x"87c0d9ff",
  1559 => x"58a6ecc0",
  1560 => x"87f8d8ff",
  1561 => x"58a6f0c0",
  1562 => x"05a8ecc0",
  1563 => x"a687c9c0",
  1564 => x"66e8c048",
  1565 => x"87c4c078",
  1566 => x"87f9d5ff",
  1567 => x"cc4966d0",
  1568 => x"66c4c191",
  1569 => x"c8807148",
  1570 => x"66c458a6",
  1571 => x"c482c84a",
  1572 => x"81ca4966",
  1573 => x"5166e8c0",
  1574 => x"4966ecc0",
  1575 => x"e8c081c1",
  1576 => x"48c18966",
  1577 => x"49703071",
  1578 => x"977189c1",
  1579 => x"e4eec27a",
  1580 => x"e8c049bf",
  1581 => x"6a972966",
  1582 => x"9871484a",
  1583 => x"58a6f4c0",
  1584 => x"c44866c4",
  1585 => x"58a6cc80",
  1586 => x"4dbf66c8",
  1587 => x"4866e0c0",
  1588 => x"c002a86e",
  1589 => x"7ec087c5",
  1590 => x"c187c2c0",
  1591 => x"c01e6e7e",
  1592 => x"49751ee0",
  1593 => x"87c9d5ff",
  1594 => x"4c7086c8",
  1595 => x"06acb7c0",
  1596 => x"7487d4c1",
  1597 => x"bf66c885",
  1598 => x"81e0c049",
  1599 => x"c14b8975",
  1600 => x"714acce9",
  1601 => x"87dce0fe",
  1602 => x"7e7585c2",
  1603 => x"4866e4c0",
  1604 => x"e8c080c1",
  1605 => x"f0c058a6",
  1606 => x"81c14966",
  1607 => x"c002a970",
  1608 => x"4dc087c5",
  1609 => x"c187c2c0",
  1610 => x"cc1e754d",
  1611 => x"c049bf66",
  1612 => x"66c481e0",
  1613 => x"c81e7189",
  1614 => x"d3ff4966",
  1615 => x"86c887f3",
  1616 => x"01a8b7c0",
  1617 => x"c087c5ff",
  1618 => x"c00266e4",
  1619 => x"66c487d3",
  1620 => x"c081c949",
  1621 => x"c45166e4",
  1622 => x"d3c14866",
  1623 => x"cec078c7",
  1624 => x"4966c487",
  1625 => x"51c281c9",
  1626 => x"c14866c4",
  1627 => x"d078c5d5",
  1628 => x"66d44866",
  1629 => x"cbc004a8",
  1630 => x"4866d087",
  1631 => x"a6d480c1",
  1632 => x"87dac058",
  1633 => x"c14866d4",
  1634 => x"58a6d888",
  1635 => x"ff87cfc0",
  1636 => x"7087cad2",
  1637 => x"87c6c04c",
  1638 => x"87c1d2ff",
  1639 => x"66dc4c70",
  1640 => x"c080c148",
  1641 => x"7458a6e0",
  1642 => x"cbc0029c",
  1643 => x"4866d087",
  1644 => x"a866ccc1",
  1645 => x"87f1f204",
  1646 => x"c74866d0",
  1647 => x"e1c003a8",
  1648 => x"4c66d087",
  1649 => x"48c8efc2",
  1650 => x"497478c0",
  1651 => x"c4c191cc",
  1652 => x"a1c48166",
  1653 => x"c04a6a4a",
  1654 => x"84c17952",
  1655 => x"ff04acc7",
  1656 => x"e0c087e2",
  1657 => x"e2c00266",
  1658 => x"66c4c187",
  1659 => x"81d4c149",
  1660 => x"4a66c4c1",
  1661 => x"c082dcc1",
  1662 => x"f9d1c152",
  1663 => x"66c4c179",
  1664 => x"81d8c149",
  1665 => x"79d0e9c1",
  1666 => x"c187d6c0",
  1667 => x"c14966c4",
  1668 => x"c4c181d4",
  1669 => x"d8c14a66",
  1670 => x"d8e9c182",
  1671 => x"f0d1c17a",
  1672 => x"d7d5c179",
  1673 => x"66c4c14a",
  1674 => x"81e0c149",
  1675 => x"cfff7972",
  1676 => x"66cc87e2",
  1677 => x"8eccff48",
  1678 => x"4c264d26",
  1679 => x"4f264b26",
  1680 => x"64616f4c",
  1681 => x"202e2a20",
  1682 => x"00000000",
  1683 => x"0000203a",
  1684 => x"61422080",
  1685 => x"00006b63",
  1686 => x"78452080",
  1687 => x"1e007469",
  1688 => x"efc21ec7",
  1689 => x"c11ebfc4",
  1690 => x"c21ee4ed",
  1691 => x"bf97e8ee",
  1692 => x"87f5ec49",
  1693 => x"49e4edc1",
  1694 => x"87dee2c0",
  1695 => x"4f268ef4",
  1696 => x"c01e731e",
  1697 => x"d8edc14b",
  1698 => x"c150c048",
  1699 => x"49bfd0ef",
  1700 => x"87f6d3ff",
  1701 => x"c4059870",
  1702 => x"e4eac187",
  1703 => x"2648734b",
  1704 => x"004f264b",
  1705 => x"204d4f52",
  1706 => x"64616f6c",
  1707 => x"20676e69",
  1708 => x"6c696166",
  1709 => x"1e006465",
  1710 => x"d0c81e73",
  1711 => x"d0efc287",
  1712 => x"c150c048",
  1713 => x"c148fcee",
  1714 => x"fe78c4ed",
  1715 => x"c049a0e8",
  1716 => x"c787c7e1",
  1717 => x"87f4df49",
  1718 => x"e1c049c1",
  1719 => x"d4ff87cf",
  1720 => x"78ffc348",
  1721 => x"87e4e2fe",
  1722 => x"cd029870",
  1723 => x"e0ecfe87",
  1724 => x"02987087",
  1725 => x"4ac187c4",
  1726 => x"4ac087c2",
  1727 => x"c8029a72",
  1728 => x"d0edc187",
  1729 => x"ded6fe49",
  1730 => x"c4efc287",
  1731 => x"c278c048",
  1732 => x"c048e8ee",
  1733 => x"c6fd4950",
  1734 => x"87e4fd87",
  1735 => x"029b4b70",
  1736 => x"efc187cb",
  1737 => x"49c75bc0",
  1738 => x"c587e1de",
  1739 => x"df49c087",
  1740 => x"d2c387fb",
  1741 => x"dce1c087",
  1742 => x"f0eec087",
  1743 => x"87f5ff87",
  1744 => x"4f264b26",
  1745 => x"746f6f42",
  1746 => x"2e676e69",
  1747 => x"00002e2e",
  1748 => x"4f204453",
  1749 => x"0000004b",
  1750 => x"00000000",
  1751 => x"00000000",
  1752 => x"00000001",
  1753 => x"0000115e",
  1754 => x"00002bdc",
  1755 => x"00000000",
  1756 => x"0000115e",
  1757 => x"00002bfa",
  1758 => x"00000000",
  1759 => x"0000115e",
  1760 => x"00002c18",
  1761 => x"00000000",
  1762 => x"0000115e",
  1763 => x"00002c36",
  1764 => x"00000000",
  1765 => x"0000115e",
  1766 => x"00002c54",
  1767 => x"00000000",
  1768 => x"0000115e",
  1769 => x"00002c72",
  1770 => x"00000000",
  1771 => x"0000115e",
  1772 => x"00002c90",
  1773 => x"00000000",
  1774 => x"00001479",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00001213",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00001bd4",
  1781 => x"20434242",
  1782 => x"20202020",
  1783 => x"004d4f52",
  1784 => x"db86fc1e",
  1785 => x"fc7e7087",
  1786 => x"1e4f268e",
  1787 => x"c048f0fe",
  1788 => x"7909cd78",
  1789 => x"1e4f2609",
  1790 => x"49e0efc1",
  1791 => x"4f2687ed",
  1792 => x"bff0fe1e",
  1793 => x"1e4f2648",
  1794 => x"c148f0fe",
  1795 => x"1e4f2678",
  1796 => x"c048f0fe",
  1797 => x"1e4f2678",
  1798 => x"52c04a71",
  1799 => x"0e4f2651",
  1800 => x"5d5c5b5e",
  1801 => x"7186f40e",
  1802 => x"7e6d974d",
  1803 => x"974ca5c1",
  1804 => x"a6c8486c",
  1805 => x"c4486e58",
  1806 => x"c505a866",
  1807 => x"c048ff87",
  1808 => x"caff87e6",
  1809 => x"49a5c287",
  1810 => x"714b6c97",
  1811 => x"6b974ba3",
  1812 => x"7e6c974b",
  1813 => x"80c1486e",
  1814 => x"c758a6c8",
  1815 => x"58a6cc98",
  1816 => x"fe7c9770",
  1817 => x"487387e1",
  1818 => x"4d268ef4",
  1819 => x"4b264c26",
  1820 => x"5e0e4f26",
  1821 => x"f40e5c5b",
  1822 => x"d84c7186",
  1823 => x"ffc34a66",
  1824 => x"4ba4c29a",
  1825 => x"73496c97",
  1826 => x"517249a1",
  1827 => x"6e7e6c97",
  1828 => x"c880c148",
  1829 => x"98c758a6",
  1830 => x"7058a6cc",
  1831 => x"268ef454",
  1832 => x"264b264c",
  1833 => x"86fc1e4f",
  1834 => x"e087e4fd",
  1835 => x"c0494abf",
  1836 => x"0299c0e0",
  1837 => x"1e7287cb",
  1838 => x"49f0f2c2",
  1839 => x"c487f3fe",
  1840 => x"87fcfc86",
  1841 => x"fefc7e70",
  1842 => x"268efc87",
  1843 => x"f2c21e4f",
  1844 => x"c2fd49f0",
  1845 => x"e5f2c187",
  1846 => x"87cffc49",
  1847 => x"2687f1c2",
  1848 => x"1e731e4f",
  1849 => x"49f0f2c2",
  1850 => x"7087f4fc",
  1851 => x"aab7c04a",
  1852 => x"87ccc204",
  1853 => x"05aaf0c3",
  1854 => x"f6c187c9",
  1855 => x"78c148c8",
  1856 => x"c387edc1",
  1857 => x"c905aae0",
  1858 => x"ccf6c187",
  1859 => x"c178c148",
  1860 => x"f6c187de",
  1861 => x"c602bfcc",
  1862 => x"a2c0c287",
  1863 => x"7287c24b",
  1864 => x"c8f6c14b",
  1865 => x"e0c002bf",
  1866 => x"c4497387",
  1867 => x"c19129b7",
  1868 => x"7381e4f7",
  1869 => x"c29acf4a",
  1870 => x"7248c192",
  1871 => x"ff4a7030",
  1872 => x"694872ba",
  1873 => x"db797098",
  1874 => x"c4497387",
  1875 => x"c19129b7",
  1876 => x"7381e4f7",
  1877 => x"c29acf4a",
  1878 => x"7248c392",
  1879 => x"484a7030",
  1880 => x"7970b069",
  1881 => x"48ccf6c1",
  1882 => x"f6c178c0",
  1883 => x"78c048c8",
  1884 => x"49f0f2c2",
  1885 => x"7087e8fa",
  1886 => x"aab7c04a",
  1887 => x"87f4fd03",
  1888 => x"4b2648c0",
  1889 => x"00004f26",
  1890 => x"00000000",
  1891 => x"00000000",
  1892 => x"724ac01e",
  1893 => x"c191c449",
  1894 => x"c081e4f7",
  1895 => x"d082c179",
  1896 => x"ee04aab7",
  1897 => x"0e4f2687",
  1898 => x"5d5c5b5e",
  1899 => x"f94d710e",
  1900 => x"4a7587dd",
  1901 => x"922ab7c4",
  1902 => x"82e4f7c1",
  1903 => x"9ccf4c75",
  1904 => x"496a94c2",
  1905 => x"c32b744b",
  1906 => x"7448c29b",
  1907 => x"ff4c7030",
  1908 => x"714874bc",
  1909 => x"f87a7098",
  1910 => x"487387ed",
  1911 => x"4c264d26",
  1912 => x"4f264b26",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"00000000",
  1926 => x"00000000",
  1927 => x"00000000",
  1928 => x"00000000",
  1929 => x"48d0ff1e",
  1930 => x"7178e1c8",
  1931 => x"08d4ff48",
  1932 => x"1e4f2678",
  1933 => x"c848d0ff",
  1934 => x"487178e1",
  1935 => x"7808d4ff",
  1936 => x"ff4866c4",
  1937 => x"267808d4",
  1938 => x"4a711e4f",
  1939 => x"1e4966c4",
  1940 => x"deff4972",
  1941 => x"48d0ff87",
  1942 => x"fc78e0c0",
  1943 => x"1e4f268e",
  1944 => x"4b711e73",
  1945 => x"1e4966c8",
  1946 => x"e0c14a73",
  1947 => x"d8ff49a2",
  1948 => x"268efc87",
  1949 => x"1e4f264b",
  1950 => x"c848d0ff",
  1951 => x"487178c9",
  1952 => x"7808d4ff",
  1953 => x"711e4f26",
  1954 => x"87eb494a",
  1955 => x"c848d0ff",
  1956 => x"1e4f2678",
  1957 => x"4b711e73",
  1958 => x"bfc8f3c2",
  1959 => x"c287c302",
  1960 => x"d0ff87eb",
  1961 => x"78c9c848",
  1962 => x"e0c04873",
  1963 => x"08d4ffb0",
  1964 => x"fcf2c278",
  1965 => x"c878c048",
  1966 => x"87c50266",
  1967 => x"c249ffc3",
  1968 => x"c249c087",
  1969 => x"cc59c4f3",
  1970 => x"87c60266",
  1971 => x"4ad5d5c5",
  1972 => x"ffcf87c4",
  1973 => x"f3c24aff",
  1974 => x"f3c25ac8",
  1975 => x"78c148c8",
  1976 => x"4f264b26",
  1977 => x"5c5b5e0e",
  1978 => x"4d710e5d",
  1979 => x"bfc4f3c2",
  1980 => x"029d754b",
  1981 => x"c84987cb",
  1982 => x"ccfac191",
  1983 => x"c482714a",
  1984 => x"ccfec187",
  1985 => x"124cc04a",
  1986 => x"c2997349",
  1987 => x"48bfc0f3",
  1988 => x"d4ffb871",
  1989 => x"b7c17808",
  1990 => x"b7c8842b",
  1991 => x"87e704ac",
  1992 => x"bffcf2c2",
  1993 => x"c280c848",
  1994 => x"2658c0f3",
  1995 => x"264c264d",
  1996 => x"1e4f264b",
  1997 => x"4b711e73",
  1998 => x"029a4a13",
  1999 => x"497287cb",
  2000 => x"1387e1fe",
  2001 => x"f5059a4a",
  2002 => x"264b2687",
  2003 => x"f2c21e4f",
  2004 => x"c249bffc",
  2005 => x"c148fcf2",
  2006 => x"c0c478a1",
  2007 => x"db03a9b7",
  2008 => x"48d4ff87",
  2009 => x"bfc0f3c2",
  2010 => x"fcf2c278",
  2011 => x"f2c249bf",
  2012 => x"a1c148fc",
  2013 => x"b7c0c478",
  2014 => x"87e504a9",
  2015 => x"c848d0ff",
  2016 => x"c8f3c278",
  2017 => x"2678c048",
  2018 => x"0000004f",
  2019 => x"00000000",
  2020 => x"00000000",
  2021 => x"5f000000",
  2022 => x"0000005f",
  2023 => x"00030300",
  2024 => x"00000303",
  2025 => x"147f7f14",
  2026 => x"00147f7f",
  2027 => x"6b2e2400",
  2028 => x"00123a6b",
  2029 => x"18366a4c",
  2030 => x"0032566c",
  2031 => x"594f7e30",
  2032 => x"40683a77",
  2033 => x"07040000",
  2034 => x"00000003",
  2035 => x"3e1c0000",
  2036 => x"00004163",
  2037 => x"63410000",
  2038 => x"00001c3e",
  2039 => x"1c3e2a08",
  2040 => x"082a3e1c",
  2041 => x"3e080800",
  2042 => x"0008083e",
  2043 => x"e0800000",
  2044 => x"00000060",
  2045 => x"08080800",
  2046 => x"00080808",
  2047 => x"60000000",
  2048 => x"00000060",
  2049 => x"18306040",
  2050 => x"0103060c",
  2051 => x"597f3e00",
  2052 => x"003e7f4d",
  2053 => x"7f060400",
  2054 => x"0000007f",
  2055 => x"71634200",
  2056 => x"00464f59",
  2057 => x"49632200",
  2058 => x"00367f49",
  2059 => x"13161c18",
  2060 => x"00107f7f",
  2061 => x"45672700",
  2062 => x"00397d45",
  2063 => x"4b7e3c00",
  2064 => x"00307949",
  2065 => x"71010100",
  2066 => x"00070f79",
  2067 => x"497f3600",
  2068 => x"00367f49",
  2069 => x"494f0600",
  2070 => x"001e3f69",
  2071 => x"66000000",
  2072 => x"00000066",
  2073 => x"e6800000",
  2074 => x"00000066",
  2075 => x"14080800",
  2076 => x"00222214",
  2077 => x"14141400",
  2078 => x"00141414",
  2079 => x"14222200",
  2080 => x"00080814",
  2081 => x"51030200",
  2082 => x"00060f59",
  2083 => x"5d417f3e",
  2084 => x"001e1f55",
  2085 => x"097f7e00",
  2086 => x"007e7f09",
  2087 => x"497f7f00",
  2088 => x"00367f49",
  2089 => x"633e1c00",
  2090 => x"00414141",
  2091 => x"417f7f00",
  2092 => x"001c3e63",
  2093 => x"497f7f00",
  2094 => x"00414149",
  2095 => x"097f7f00",
  2096 => x"00010109",
  2097 => x"417f3e00",
  2098 => x"007a7b49",
  2099 => x"087f7f00",
  2100 => x"007f7f08",
  2101 => x"7f410000",
  2102 => x"0000417f",
  2103 => x"40602000",
  2104 => x"003f7f40",
  2105 => x"1c087f7f",
  2106 => x"00416336",
  2107 => x"407f7f00",
  2108 => x"00404040",
  2109 => x"0c067f7f",
  2110 => x"007f7f06",
  2111 => x"0c067f7f",
  2112 => x"007f7f18",
  2113 => x"417f3e00",
  2114 => x"003e7f41",
  2115 => x"097f7f00",
  2116 => x"00060f09",
  2117 => x"61417f3e",
  2118 => x"00407e7f",
  2119 => x"097f7f00",
  2120 => x"00667f19",
  2121 => x"4d6f2600",
  2122 => x"00327b59",
  2123 => x"7f010100",
  2124 => x"0001017f",
  2125 => x"407f3f00",
  2126 => x"003f7f40",
  2127 => x"703f0f00",
  2128 => x"000f3f70",
  2129 => x"18307f7f",
  2130 => x"007f7f30",
  2131 => x"1c366341",
  2132 => x"4163361c",
  2133 => x"7c060301",
  2134 => x"0103067c",
  2135 => x"4d597161",
  2136 => x"00414347",
  2137 => x"7f7f0000",
  2138 => x"00004141",
  2139 => x"0c060301",
  2140 => x"40603018",
  2141 => x"41410000",
  2142 => x"00007f7f",
  2143 => x"03060c08",
  2144 => x"00080c06",
  2145 => x"80808080",
  2146 => x"00808080",
  2147 => x"03000000",
  2148 => x"00000407",
  2149 => x"54742000",
  2150 => x"00787c54",
  2151 => x"447f7f00",
  2152 => x"00387c44",
  2153 => x"447c3800",
  2154 => x"00004444",
  2155 => x"447c3800",
  2156 => x"007f7f44",
  2157 => x"547c3800",
  2158 => x"00185c54",
  2159 => x"7f7e0400",
  2160 => x"00000505",
  2161 => x"a4bc1800",
  2162 => x"007cfca4",
  2163 => x"047f7f00",
  2164 => x"00787c04",
  2165 => x"3d000000",
  2166 => x"0000407d",
  2167 => x"80808000",
  2168 => x"00007dfd",
  2169 => x"107f7f00",
  2170 => x"00446c38",
  2171 => x"3f000000",
  2172 => x"0000407f",
  2173 => x"180c7c7c",
  2174 => x"00787c0c",
  2175 => x"047c7c00",
  2176 => x"00787c04",
  2177 => x"447c3800",
  2178 => x"00387c44",
  2179 => x"24fcfc00",
  2180 => x"00183c24",
  2181 => x"243c1800",
  2182 => x"00fcfc24",
  2183 => x"047c7c00",
  2184 => x"00080c04",
  2185 => x"545c4800",
  2186 => x"00207454",
  2187 => x"7f3f0400",
  2188 => x"00004444",
  2189 => x"407c3c00",
  2190 => x"007c7c40",
  2191 => x"603c1c00",
  2192 => x"001c3c60",
  2193 => x"30607c3c",
  2194 => x"003c7c60",
  2195 => x"10386c44",
  2196 => x"00446c38",
  2197 => x"e0bc1c00",
  2198 => x"001c3c60",
  2199 => x"74644400",
  2200 => x"00444c5c",
  2201 => x"3e080800",
  2202 => x"00414177",
  2203 => x"7f000000",
  2204 => x"0000007f",
  2205 => x"77414100",
  2206 => x"0008083e",
  2207 => x"03010102",
  2208 => x"00010202",
  2209 => x"7f7f7f7f",
  2210 => x"007f7f7f",
  2211 => x"1c1c0808",
  2212 => x"7f7f3e3e",
  2213 => x"3e3e7f7f",
  2214 => x"08081c1c",
  2215 => x"7c181000",
  2216 => x"0010187c",
  2217 => x"7c301000",
  2218 => x"0010307c",
  2219 => x"60603010",
  2220 => x"00061e78",
  2221 => x"183c6642",
  2222 => x"0042663c",
  2223 => x"c26a3878",
  2224 => x"00386cc6",
  2225 => x"60000060",
  2226 => x"00600000",
  2227 => x"5c5b5e0e",
  2228 => x"86fc0e5d",
  2229 => x"f3c27e71",
  2230 => x"c04cbfd0",
  2231 => x"c41ec04b",
  2232 => x"c402ab66",
  2233 => x"c24dc087",
  2234 => x"754dc187",
  2235 => x"ee49731e",
  2236 => x"86c887e1",
  2237 => x"ef49e0c0",
  2238 => x"a4c487ea",
  2239 => x"f0496a4a",
  2240 => x"c8f187f1",
  2241 => x"c184cc87",
  2242 => x"abb7c883",
  2243 => x"87cdff04",
  2244 => x"4d268efc",
  2245 => x"4b264c26",
  2246 => x"711e4f26",
  2247 => x"d4f3c24a",
  2248 => x"d4f3c25a",
  2249 => x"4978c748",
  2250 => x"2687e1fe",
  2251 => x"1e731e4f",
  2252 => x"b7c04a71",
  2253 => x"87d303aa",
  2254 => x"bfd0d9c2",
  2255 => x"c187c405",
  2256 => x"c087c24b",
  2257 => x"d4d9c24b",
  2258 => x"c287c45b",
  2259 => x"fc5ad4d9",
  2260 => x"d0d9c248",
  2261 => x"c14a78bf",
  2262 => x"a2c0c19a",
  2263 => x"87e6ec49",
  2264 => x"4f264b26",
  2265 => x"c44a711e",
  2266 => x"49721e66",
  2267 => x"fc87f0eb",
  2268 => x"1e4f268e",
  2269 => x"c348d4ff",
  2270 => x"d0ff78ff",
  2271 => x"78e1c048",
  2272 => x"c148d4ff",
  2273 => x"c4487178",
  2274 => x"08d4ff30",
  2275 => x"48d0ff78",
  2276 => x"2678e0c0",
  2277 => x"5b5e0e4f",
  2278 => x"f00e5d5c",
  2279 => x"48a6c886",
  2280 => x"ec4d78c0",
  2281 => x"80fc7ebf",
  2282 => x"bfd0f3c2",
  2283 => x"4cbfe878",
  2284 => x"bfd0d9c2",
  2285 => x"87e9e449",
  2286 => x"ca49eecb",
  2287 => x"4b7087d6",
  2288 => x"e2e749c7",
  2289 => x"05987087",
  2290 => x"496e87c8",
  2291 => x"c10299c1",
  2292 => x"4dc187c1",
  2293 => x"c27ebfec",
  2294 => x"49bfd0d9",
  2295 => x"7387c2e4",
  2296 => x"87fcc949",
  2297 => x"d7029870",
  2298 => x"c8d9c287",
  2299 => x"b9c149bf",
  2300 => x"59ccd9c2",
  2301 => x"87fbfd71",
  2302 => x"c949eecb",
  2303 => x"4b7087d6",
  2304 => x"e2e649c7",
  2305 => x"05987087",
  2306 => x"6e87c7ff",
  2307 => x"0599c149",
  2308 => x"7587fffe",
  2309 => x"e3c0029d",
  2310 => x"d0d9c287",
  2311 => x"bac14abf",
  2312 => x"5ad4d9c2",
  2313 => x"0a7a0afc",
  2314 => x"c0c19ac1",
  2315 => x"d5e949a2",
  2316 => x"49dac187",
  2317 => x"c887f0e5",
  2318 => x"78c148a6",
  2319 => x"bfd0d9c2",
  2320 => x"87e9c005",
  2321 => x"ffc34974",
  2322 => x"c01e7199",
  2323 => x"87d4fc49",
  2324 => x"b7c84974",
  2325 => x"c11e7129",
  2326 => x"87c8fc49",
  2327 => x"fdc386c8",
  2328 => x"87c3e549",
  2329 => x"e449fac3",
  2330 => x"d1c787fd",
  2331 => x"c3497487",
  2332 => x"b7c899ff",
  2333 => x"74b4712c",
  2334 => x"87df029c",
  2335 => x"bfccd9c2",
  2336 => x"87dcc749",
  2337 => x"c0059870",
  2338 => x"4cc087c4",
  2339 => x"e0c287d3",
  2340 => x"87c0c749",
  2341 => x"58d0d9c2",
  2342 => x"c287c6c0",
  2343 => x"c048ccd9",
  2344 => x"c8497478",
  2345 => x"87ce0599",
  2346 => x"e349f5c3",
  2347 => x"497087f9",
  2348 => x"c00299c2",
  2349 => x"f3c287e9",
  2350 => x"c002bfd4",
  2351 => x"c14887c9",
  2352 => x"d8f3c288",
  2353 => x"c487d358",
  2354 => x"e0c14866",
  2355 => x"6e7e7080",
  2356 => x"c5c002bf",
  2357 => x"49ff4b87",
  2358 => x"a6c80f73",
  2359 => x"7478c148",
  2360 => x"0599c449",
  2361 => x"c387cec0",
  2362 => x"fae249f2",
  2363 => x"c2497087",
  2364 => x"f0c00299",
  2365 => x"d4f3c287",
  2366 => x"c7487ebf",
  2367 => x"c003a8b7",
  2368 => x"486e87cb",
  2369 => x"f3c280c1",
  2370 => x"d3c058d8",
  2371 => x"4866c487",
  2372 => x"7080e0c1",
  2373 => x"02bf6e7e",
  2374 => x"4b87c5c0",
  2375 => x"0f7349fe",
  2376 => x"c148a6c8",
  2377 => x"49fdc378",
  2378 => x"7087fce1",
  2379 => x"0299c249",
  2380 => x"c287e9c0",
  2381 => x"02bfd4f3",
  2382 => x"c287c9c0",
  2383 => x"c048d4f3",
  2384 => x"87d3c078",
  2385 => x"c14866c4",
  2386 => x"7e7080e0",
  2387 => x"c002bf6e",
  2388 => x"fd4b87c5",
  2389 => x"c80f7349",
  2390 => x"78c148a6",
  2391 => x"e149fac3",
  2392 => x"497087c5",
  2393 => x"c00299c2",
  2394 => x"f3c287ea",
  2395 => x"c748bfd4",
  2396 => x"c003a8b7",
  2397 => x"f3c287c9",
  2398 => x"78c748d4",
  2399 => x"c487d0c0",
  2400 => x"e0c14a66",
  2401 => x"c0026a82",
  2402 => x"fc4b87c5",
  2403 => x"c80f7349",
  2404 => x"78c148a6",
  2405 => x"f3c24dc0",
  2406 => x"50c048cc",
  2407 => x"c249eecb",
  2408 => x"4b7087f2",
  2409 => x"97ccf3c2",
  2410 => x"ddc105bf",
  2411 => x"c3497487",
  2412 => x"c00599f0",
  2413 => x"dac187cd",
  2414 => x"eadfff49",
  2415 => x"02987087",
  2416 => x"c187c7c1",
  2417 => x"4cbfe84d",
  2418 => x"99ffc349",
  2419 => x"712cb7c8",
  2420 => x"d0d9c2b4",
  2421 => x"dcff49bf",
  2422 => x"497387c7",
  2423 => x"7087c1c2",
  2424 => x"c6c00298",
  2425 => x"ccf3c287",
  2426 => x"c250c148",
  2427 => x"bf97ccf3",
  2428 => x"87d6c005",
  2429 => x"f0c34974",
  2430 => x"c6ff0599",
  2431 => x"49dac187",
  2432 => x"87e3deff",
  2433 => x"fe059870",
  2434 => x"9d7587f9",
  2435 => x"87e0c002",
  2436 => x"c248a6cc",
  2437 => x"78bfd4f3",
  2438 => x"cc4966cc",
  2439 => x"4866c491",
  2440 => x"7e708071",
  2441 => x"c002bf6e",
  2442 => x"cc4b87c6",
  2443 => x"0f734966",
  2444 => x"c00266c8",
  2445 => x"f3c287c8",
  2446 => x"f249bfd4",
  2447 => x"8ef087ce",
  2448 => x"4c264d26",
  2449 => x"4f264b26",
  2450 => x"00000000",
  2451 => x"00000000",
  2452 => x"00000000",
  2453 => x"ff4a711e",
  2454 => x"7249bfc8",
  2455 => x"4f2648a1",
  2456 => x"bfc8ff1e",
  2457 => x"c0c0fe89",
  2458 => x"a9c0c0c0",
  2459 => x"c087c401",
  2460 => x"c187c24a",
  2461 => x"2648724a",
  2462 => x"5b5e0e4f",
  2463 => x"710e5d5c",
  2464 => x"4cd4ff4b",
  2465 => x"c04866d0",
  2466 => x"ff49d678",
  2467 => x"c387d5de",
  2468 => x"496c7cff",
  2469 => x"7199ffc3",
  2470 => x"f0c3494d",
  2471 => x"a9e0c199",
  2472 => x"c387cb05",
  2473 => x"486c7cff",
  2474 => x"66d098c3",
  2475 => x"ffc37808",
  2476 => x"494a6c7c",
  2477 => x"ffc331c8",
  2478 => x"714a6c7c",
  2479 => x"c84972b2",
  2480 => x"7cffc331",
  2481 => x"b2714a6c",
  2482 => x"31c84972",
  2483 => x"6c7cffc3",
  2484 => x"ffb2714a",
  2485 => x"e0c048d0",
  2486 => x"029b7378",
  2487 => x"7b7287c2",
  2488 => x"4d264875",
  2489 => x"4b264c26",
  2490 => x"261e4f26",
  2491 => x"5b5e0e4f",
  2492 => x"86f80e5c",
  2493 => x"a6c81e76",
  2494 => x"87fdfd49",
  2495 => x"4b7086c4",
  2496 => x"a8c2486e",
  2497 => x"87f0c203",
  2498 => x"f0c34a73",
  2499 => x"aad0c19a",
  2500 => x"c187c702",
  2501 => x"c205aae0",
  2502 => x"497387de",
  2503 => x"c30299c8",
  2504 => x"87c6ff87",
  2505 => x"9cc34c73",
  2506 => x"c105acc2",
  2507 => x"66c487c2",
  2508 => x"7131c949",
  2509 => x"4a66c41e",
  2510 => x"f3c292d4",
  2511 => x"817249d8",
  2512 => x"87d5cefe",
  2513 => x"dbff49d8",
  2514 => x"c0c887da",
  2515 => x"f0e1c21e",
  2516 => x"c2e8fd49",
  2517 => x"48d0ff87",
  2518 => x"c278e0c0",
  2519 => x"cc1ef0e1",
  2520 => x"92d44a66",
  2521 => x"49d8f3c2",
  2522 => x"ccfe8172",
  2523 => x"86cc87dc",
  2524 => x"c105acc1",
  2525 => x"66c487c2",
  2526 => x"7131c949",
  2527 => x"4a66c41e",
  2528 => x"f3c292d4",
  2529 => x"817249d8",
  2530 => x"87cdcdfe",
  2531 => x"1ef0e1c2",
  2532 => x"d44a66c8",
  2533 => x"d8f3c292",
  2534 => x"fe817249",
  2535 => x"d787dcca",
  2536 => x"ffd9ff49",
  2537 => x"1ec0c887",
  2538 => x"49f0e1c2",
  2539 => x"87c4e6fd",
  2540 => x"d0ff86cc",
  2541 => x"78e0c048",
  2542 => x"4c268ef8",
  2543 => x"4f264b26",
  2544 => x"5c5b5e0e",
  2545 => x"86fc0e5d",
  2546 => x"d4ff4d71",
  2547 => x"7e66d44c",
  2548 => x"a8b7c348",
  2549 => x"87e2c101",
  2550 => x"66c41e75",
  2551 => x"c293d44b",
  2552 => x"7383d8f3",
  2553 => x"ccc4fe49",
  2554 => x"49a3c887",
  2555 => x"d0ff4969",
  2556 => x"78e1c848",
  2557 => x"48717cdd",
  2558 => x"7098ffc3",
  2559 => x"c84a717c",
  2560 => x"48722ab7",
  2561 => x"7098ffc3",
  2562 => x"d04a717c",
  2563 => x"48722ab7",
  2564 => x"7098ffc3",
  2565 => x"d848717c",
  2566 => x"7c7028b7",
  2567 => x"7c7c7cc0",
  2568 => x"7c7c7c7c",
  2569 => x"7c7c7c7c",
  2570 => x"48d0ff7c",
  2571 => x"c478e0c0",
  2572 => x"49dc1e66",
  2573 => x"87d1d8ff",
  2574 => x"8efc86c8",
  2575 => x"4c264d26",
  2576 => x"4f264b26",
  2577 => x"00001bf7",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
