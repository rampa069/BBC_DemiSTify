
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"7c",x"40",x"40",x"7c"),
     1 => (x"1c",x"00",x"00",x"7c"),
     2 => (x"3c",x"60",x"60",x"3c"),
     3 => (x"7c",x"3c",x"00",x"1c"),
     4 => (x"7c",x"60",x"30",x"60"),
     5 => (x"6c",x"44",x"00",x"3c"),
     6 => (x"6c",x"38",x"10",x"38"),
     7 => (x"1c",x"00",x"00",x"44"),
     8 => (x"3c",x"60",x"e0",x"bc"),
     9 => (x"44",x"00",x"00",x"1c"),
    10 => (x"4c",x"5c",x"74",x"64"),
    11 => (x"08",x"00",x"00",x"44"),
    12 => (x"41",x"77",x"3e",x"08"),
    13 => (x"00",x"00",x"00",x"41"),
    14 => (x"00",x"7f",x"7f",x"00"),
    15 => (x"41",x"00",x"00",x"00"),
    16 => (x"08",x"3e",x"77",x"41"),
    17 => (x"01",x"02",x"00",x"08"),
    18 => (x"02",x"02",x"03",x"01"),
    19 => (x"7f",x"7f",x"00",x"01"),
    20 => (x"7f",x"7f",x"7f",x"7f"),
    21 => (x"08",x"08",x"00",x"7f"),
    22 => (x"3e",x"3e",x"1c",x"1c"),
    23 => (x"7f",x"7f",x"7f",x"7f"),
    24 => (x"1c",x"1c",x"3e",x"3e"),
    25 => (x"10",x"00",x"08",x"08"),
    26 => (x"18",x"7c",x"7c",x"18"),
    27 => (x"10",x"00",x"00",x"10"),
    28 => (x"30",x"7c",x"7c",x"30"),
    29 => (x"30",x"10",x"00",x"10"),
    30 => (x"1e",x"78",x"60",x"60"),
    31 => (x"66",x"42",x"00",x"06"),
    32 => (x"66",x"3c",x"18",x"3c"),
    33 => (x"38",x"78",x"00",x"42"),
    34 => (x"6c",x"c6",x"c2",x"6a"),
    35 => (x"00",x"60",x"00",x"38"),
    36 => (x"00",x"00",x"60",x"00"),
    37 => (x"5e",x"0e",x"00",x"60"),
    38 => (x"0e",x"5d",x"5c",x"5b"),
    39 => (x"c2",x"4c",x"71",x"1e"),
    40 => (x"4d",x"bf",x"d9",x"ee"),
    41 => (x"1e",x"c0",x"4b",x"c0"),
    42 => (x"c7",x"02",x"ab",x"74"),
    43 => (x"48",x"a6",x"c4",x"87"),
    44 => (x"87",x"c5",x"78",x"c0"),
    45 => (x"c1",x"48",x"a6",x"c4"),
    46 => (x"1e",x"66",x"c4",x"78"),
    47 => (x"df",x"ee",x"49",x"73"),
    48 => (x"c0",x"86",x"c8",x"87"),
    49 => (x"ee",x"ef",x"49",x"e0"),
    50 => (x"4a",x"a5",x"c4",x"87"),
    51 => (x"f0",x"f0",x"49",x"6a"),
    52 => (x"87",x"c6",x"f1",x"87"),
    53 => (x"83",x"c1",x"85",x"cb"),
    54 => (x"04",x"ab",x"b7",x"c8"),
    55 => (x"26",x"87",x"c7",x"ff"),
    56 => (x"4c",x"26",x"4d",x"26"),
    57 => (x"4f",x"26",x"4b",x"26"),
    58 => (x"c2",x"4a",x"71",x"1e"),
    59 => (x"c2",x"5a",x"dd",x"ee"),
    60 => (x"c7",x"48",x"dd",x"ee"),
    61 => (x"dd",x"fe",x"49",x"78"),
    62 => (x"1e",x"4f",x"26",x"87"),
    63 => (x"4a",x"71",x"1e",x"73"),
    64 => (x"03",x"aa",x"b7",x"c0"),
    65 => (x"d2",x"c2",x"87",x"d3"),
    66 => (x"c4",x"05",x"bf",x"fe"),
    67 => (x"c2",x"4b",x"c1",x"87"),
    68 => (x"c2",x"4b",x"c0",x"87"),
    69 => (x"c4",x"5b",x"c2",x"d3"),
    70 => (x"c2",x"d3",x"c2",x"87"),
    71 => (x"fe",x"d2",x"c2",x"5a"),
    72 => (x"9a",x"c1",x"4a",x"bf"),
    73 => (x"49",x"a2",x"c0",x"c1"),
    74 => (x"fc",x"87",x"e8",x"ec"),
    75 => (x"fe",x"d2",x"c2",x"48"),
    76 => (x"ef",x"fe",x"78",x"bf"),
    77 => (x"4a",x"71",x"1e",x"87"),
    78 => (x"72",x"1e",x"66",x"c4"),
    79 => (x"87",x"f9",x"ea",x"49"),
    80 => (x"1e",x"4f",x"26",x"26"),
    81 => (x"c3",x"48",x"d4",x"ff"),
    82 => (x"d0",x"ff",x"78",x"ff"),
    83 => (x"78",x"e1",x"c0",x"48"),
    84 => (x"c1",x"48",x"d4",x"ff"),
    85 => (x"c4",x"48",x"71",x"78"),
    86 => (x"08",x"d4",x"ff",x"30"),
    87 => (x"48",x"d0",x"ff",x"78"),
    88 => (x"26",x"78",x"e0",x"c0"),
    89 => (x"d2",x"c2",x"1e",x"4f"),
    90 => (x"e6",x"49",x"bf",x"fe"),
    91 => (x"ee",x"c2",x"87",x"f9"),
    92 => (x"bf",x"e8",x"48",x"d1"),
    93 => (x"cd",x"ee",x"c2",x"78"),
    94 => (x"78",x"bf",x"ec",x"48"),
    95 => (x"bf",x"d1",x"ee",x"c2"),
    96 => (x"ff",x"c3",x"49",x"4a"),
    97 => (x"2a",x"b7",x"c8",x"99"),
    98 => (x"b0",x"71",x"48",x"72"),
    99 => (x"58",x"d9",x"ee",x"c2"),
   100 => (x"5e",x"0e",x"4f",x"26"),
   101 => (x"0e",x"5d",x"5c",x"5b"),
   102 => (x"c8",x"ff",x"4b",x"71"),
   103 => (x"cc",x"ee",x"c2",x"87"),
   104 => (x"73",x"50",x"c0",x"48"),
   105 => (x"87",x"df",x"e6",x"49"),
   106 => (x"c2",x"4c",x"49",x"70"),
   107 => (x"49",x"ee",x"cb",x"9c"),
   108 => (x"70",x"87",x"d3",x"cc"),
   109 => (x"cc",x"ee",x"c2",x"4d"),
   110 => (x"c1",x"05",x"bf",x"97"),
   111 => (x"66",x"d0",x"87",x"e2"),
   112 => (x"d5",x"ee",x"c2",x"49"),
   113 => (x"d6",x"05",x"99",x"bf"),
   114 => (x"49",x"66",x"d4",x"87"),
   115 => (x"bf",x"cd",x"ee",x"c2"),
   116 => (x"87",x"cb",x"05",x"99"),
   117 => (x"ee",x"e5",x"49",x"73"),
   118 => (x"02",x"98",x"70",x"87"),
   119 => (x"c1",x"87",x"c1",x"c1"),
   120 => (x"87",x"c1",x"fe",x"4c"),
   121 => (x"e9",x"cb",x"49",x"75"),
   122 => (x"02",x"98",x"70",x"87"),
   123 => (x"ee",x"c2",x"87",x"c6"),
   124 => (x"50",x"c1",x"48",x"cc"),
   125 => (x"97",x"cc",x"ee",x"c2"),
   126 => (x"e3",x"c0",x"05",x"bf"),
   127 => (x"d5",x"ee",x"c2",x"87"),
   128 => (x"66",x"d0",x"49",x"bf"),
   129 => (x"d6",x"ff",x"05",x"99"),
   130 => (x"cd",x"ee",x"c2",x"87"),
   131 => (x"66",x"d4",x"49",x"bf"),
   132 => (x"ca",x"ff",x"05",x"99"),
   133 => (x"e4",x"49",x"73",x"87"),
   134 => (x"98",x"70",x"87",x"ed"),
   135 => (x"87",x"ff",x"fe",x"05"),
   136 => (x"fb",x"fa",x"48",x"74"),
   137 => (x"5b",x"5e",x"0e",x"87"),
   138 => (x"f8",x"0e",x"5d",x"5c"),
   139 => (x"4c",x"4d",x"c0",x"86"),
   140 => (x"c4",x"7e",x"bf",x"ec"),
   141 => (x"ee",x"c2",x"48",x"a6"),
   142 => (x"c1",x"78",x"bf",x"d9"),
   143 => (x"c7",x"1e",x"c0",x"1e"),
   144 => (x"87",x"ce",x"fd",x"49"),
   145 => (x"98",x"70",x"86",x"c8"),
   146 => (x"ff",x"87",x"cd",x"02"),
   147 => (x"87",x"eb",x"fa",x"49"),
   148 => (x"e3",x"49",x"da",x"c1"),
   149 => (x"4d",x"c1",x"87",x"f1"),
   150 => (x"97",x"cc",x"ee",x"c2"),
   151 => (x"87",x"cf",x"02",x"bf"),
   152 => (x"bf",x"e6",x"d2",x"c2"),
   153 => (x"c2",x"b9",x"c1",x"49"),
   154 => (x"71",x"59",x"ea",x"d2"),
   155 => (x"c2",x"87",x"d4",x"fb"),
   156 => (x"4b",x"bf",x"d1",x"ee"),
   157 => (x"bf",x"fe",x"d2",x"c2"),
   158 => (x"87",x"d9",x"c1",x"05"),
   159 => (x"c8",x"48",x"a6",x"c4"),
   160 => (x"c2",x"78",x"c0",x"c0"),
   161 => (x"6e",x"7e",x"ea",x"d2"),
   162 => (x"6e",x"49",x"bf",x"97"),
   163 => (x"70",x"80",x"c1",x"48"),
   164 => (x"f2",x"e2",x"71",x"7e"),
   165 => (x"02",x"98",x"70",x"87"),
   166 => (x"66",x"c4",x"87",x"c3"),
   167 => (x"48",x"66",x"c4",x"b3"),
   168 => (x"c8",x"28",x"b7",x"c1"),
   169 => (x"98",x"70",x"58",x"a6"),
   170 => (x"87",x"db",x"ff",x"05"),
   171 => (x"e2",x"49",x"fd",x"c3"),
   172 => (x"fa",x"c3",x"87",x"d5"),
   173 => (x"87",x"cf",x"e2",x"49"),
   174 => (x"ff",x"c3",x"49",x"73"),
   175 => (x"c0",x"1e",x"71",x"99"),
   176 => (x"87",x"f1",x"f9",x"49"),
   177 => (x"b7",x"c8",x"49",x"73"),
   178 => (x"c1",x"1e",x"71",x"29"),
   179 => (x"87",x"e5",x"f9",x"49"),
   180 => (x"fa",x"c5",x"86",x"c8"),
   181 => (x"d5",x"ee",x"c2",x"87"),
   182 => (x"02",x"9b",x"4b",x"bf"),
   183 => (x"d2",x"c2",x"87",x"dd"),
   184 => (x"c7",x"49",x"bf",x"fa"),
   185 => (x"98",x"70",x"87",x"ec"),
   186 => (x"c0",x"87",x"c4",x"05"),
   187 => (x"c2",x"87",x"d2",x"4b"),
   188 => (x"d1",x"c7",x"49",x"e0"),
   189 => (x"fe",x"d2",x"c2",x"87"),
   190 => (x"c2",x"87",x"c6",x"58"),
   191 => (x"c0",x"48",x"fa",x"d2"),
   192 => (x"c2",x"49",x"73",x"78"),
   193 => (x"87",x"ce",x"05",x"99"),
   194 => (x"e0",x"49",x"eb",x"c3"),
   195 => (x"49",x"70",x"87",x"f9"),
   196 => (x"c0",x"02",x"99",x"c2"),
   197 => (x"4c",x"fb",x"87",x"c2"),
   198 => (x"99",x"c1",x"49",x"73"),
   199 => (x"c3",x"87",x"ce",x"05"),
   200 => (x"e2",x"e0",x"49",x"f4"),
   201 => (x"c2",x"49",x"70",x"87"),
   202 => (x"c2",x"c0",x"02",x"99"),
   203 => (x"73",x"4c",x"fa",x"87"),
   204 => (x"05",x"99",x"c8",x"49"),
   205 => (x"f5",x"c3",x"87",x"cd"),
   206 => (x"87",x"cb",x"e0",x"49"),
   207 => (x"99",x"c2",x"49",x"70"),
   208 => (x"c2",x"87",x"d6",x"02"),
   209 => (x"02",x"bf",x"dd",x"ee"),
   210 => (x"48",x"87",x"ca",x"c0"),
   211 => (x"ee",x"c2",x"88",x"c1"),
   212 => (x"c2",x"c0",x"58",x"e1"),
   213 => (x"c1",x"4c",x"ff",x"87"),
   214 => (x"c4",x"49",x"73",x"4d"),
   215 => (x"ce",x"c0",x"05",x"99"),
   216 => (x"49",x"f2",x"c3",x"87"),
   217 => (x"87",x"df",x"df",x"ff"),
   218 => (x"99",x"c2",x"49",x"70"),
   219 => (x"c2",x"87",x"dc",x"02"),
   220 => (x"7e",x"bf",x"dd",x"ee"),
   221 => (x"a8",x"b7",x"c7",x"48"),
   222 => (x"87",x"cb",x"c0",x"03"),
   223 => (x"80",x"c1",x"48",x"6e"),
   224 => (x"58",x"e1",x"ee",x"c2"),
   225 => (x"fe",x"87",x"c2",x"c0"),
   226 => (x"c3",x"4d",x"c1",x"4c"),
   227 => (x"de",x"ff",x"49",x"fd"),
   228 => (x"49",x"70",x"87",x"f5"),
   229 => (x"c0",x"02",x"99",x"c2"),
   230 => (x"ee",x"c2",x"87",x"d5"),
   231 => (x"c0",x"02",x"bf",x"dd"),
   232 => (x"ee",x"c2",x"87",x"c9"),
   233 => (x"78",x"c0",x"48",x"dd"),
   234 => (x"fd",x"87",x"c2",x"c0"),
   235 => (x"c3",x"4d",x"c1",x"4c"),
   236 => (x"de",x"ff",x"49",x"fa"),
   237 => (x"49",x"70",x"87",x"d1"),
   238 => (x"c0",x"02",x"99",x"c2"),
   239 => (x"ee",x"c2",x"87",x"d9"),
   240 => (x"c7",x"48",x"bf",x"dd"),
   241 => (x"c0",x"03",x"a8",x"b7"),
   242 => (x"ee",x"c2",x"87",x"c9"),
   243 => (x"78",x"c7",x"48",x"dd"),
   244 => (x"fc",x"87",x"c2",x"c0"),
   245 => (x"c0",x"4d",x"c1",x"4c"),
   246 => (x"c0",x"03",x"ac",x"b7"),
   247 => (x"66",x"c4",x"87",x"d3"),
   248 => (x"80",x"d8",x"c1",x"48"),
   249 => (x"bf",x"6e",x"7e",x"70"),
   250 => (x"87",x"c5",x"c0",x"02"),
   251 => (x"73",x"49",x"74",x"4b"),
   252 => (x"c3",x"1e",x"c0",x"0f"),
   253 => (x"da",x"c1",x"1e",x"f0"),
   254 => (x"87",x"d6",x"f6",x"49"),
   255 => (x"98",x"70",x"86",x"c8"),
   256 => (x"87",x"d8",x"c0",x"02"),
   257 => (x"bf",x"dd",x"ee",x"c2"),
   258 => (x"cb",x"49",x"6e",x"7e"),
   259 => (x"4a",x"66",x"c4",x"91"),
   260 => (x"02",x"6a",x"82",x"71"),
   261 => (x"4b",x"87",x"c5",x"c0"),
   262 => (x"0f",x"73",x"49",x"6e"),
   263 => (x"c0",x"02",x"9d",x"75"),
   264 => (x"ee",x"c2",x"87",x"c8"),
   265 => (x"f1",x"49",x"bf",x"dd"),
   266 => (x"d3",x"c2",x"87",x"ec"),
   267 => (x"c0",x"02",x"bf",x"c2"),
   268 => (x"c2",x"49",x"87",x"dd"),
   269 => (x"98",x"70",x"87",x"dc"),
   270 => (x"87",x"d3",x"c0",x"02"),
   271 => (x"bf",x"dd",x"ee",x"c2"),
   272 => (x"87",x"d2",x"f1",x"49"),
   273 => (x"f2",x"f2",x"49",x"c0"),
   274 => (x"c2",x"d3",x"c2",x"87"),
   275 => (x"f8",x"78",x"c0",x"48"),
   276 => (x"87",x"cc",x"f2",x"8e"),
   277 => (x"5c",x"5b",x"5e",x"0e"),
   278 => (x"71",x"1e",x"0e",x"5d"),
   279 => (x"d9",x"ee",x"c2",x"4c"),
   280 => (x"cd",x"c1",x"49",x"bf"),
   281 => (x"d1",x"c1",x"4d",x"a1"),
   282 => (x"74",x"7e",x"69",x"81"),
   283 => (x"87",x"cf",x"02",x"9c"),
   284 => (x"74",x"4b",x"a5",x"c4"),
   285 => (x"d9",x"ee",x"c2",x"7b"),
   286 => (x"eb",x"f1",x"49",x"bf"),
   287 => (x"74",x"7b",x"6e",x"87"),
   288 => (x"87",x"c4",x"05",x"9c"),
   289 => (x"87",x"c2",x"4b",x"c0"),
   290 => (x"49",x"73",x"4b",x"c1"),
   291 => (x"d4",x"87",x"ec",x"f1"),
   292 => (x"87",x"c8",x"02",x"66"),
   293 => (x"87",x"ee",x"c0",x"49"),
   294 => (x"87",x"c2",x"4a",x"70"),
   295 => (x"d3",x"c2",x"4a",x"c0"),
   296 => (x"f0",x"26",x"5a",x"c6"),
   297 => (x"00",x"00",x"87",x"fa"),
   298 => (x"12",x"58",x"00",x"00"),
   299 => (x"1b",x"1d",x"14",x"11"),
   300 => (x"59",x"5a",x"23",x"1c"),
   301 => (x"f2",x"f5",x"94",x"91"),
   302 => (x"00",x"00",x"f4",x"eb"),
   303 => (x"00",x"00",x"00",x"00"),
   304 => (x"00",x"00",x"00",x"00"),
   305 => (x"71",x"1e",x"00",x"00"),
   306 => (x"bf",x"c8",x"ff",x"4a"),
   307 => (x"48",x"a1",x"72",x"49"),
   308 => (x"ff",x"1e",x"4f",x"26"),
   309 => (x"fe",x"89",x"bf",x"c8"),
   310 => (x"c0",x"c0",x"c0",x"c0"),
   311 => (x"c4",x"01",x"a9",x"c0"),
   312 => (x"c2",x"4a",x"c0",x"87"),
   313 => (x"72",x"4a",x"c1",x"87"),
   314 => (x"0e",x"4f",x"26",x"48"),
   315 => (x"5d",x"5c",x"5b",x"5e"),
   316 => (x"ff",x"4b",x"71",x"0e"),
   317 => (x"66",x"d0",x"4c",x"d4"),
   318 => (x"d6",x"78",x"c0",x"48"),
   319 => (x"fe",x"da",x"ff",x"49"),
   320 => (x"7c",x"ff",x"c3",x"87"),
   321 => (x"ff",x"c3",x"49",x"6c"),
   322 => (x"49",x"4d",x"71",x"99"),
   323 => (x"c1",x"99",x"f0",x"c3"),
   324 => (x"cb",x"05",x"a9",x"e0"),
   325 => (x"7c",x"ff",x"c3",x"87"),
   326 => (x"98",x"c3",x"48",x"6c"),
   327 => (x"78",x"08",x"66",x"d0"),
   328 => (x"6c",x"7c",x"ff",x"c3"),
   329 => (x"31",x"c8",x"49",x"4a"),
   330 => (x"6c",x"7c",x"ff",x"c3"),
   331 => (x"72",x"b2",x"71",x"4a"),
   332 => (x"c3",x"31",x"c8",x"49"),
   333 => (x"4a",x"6c",x"7c",x"ff"),
   334 => (x"49",x"72",x"b2",x"71"),
   335 => (x"ff",x"c3",x"31",x"c8"),
   336 => (x"71",x"4a",x"6c",x"7c"),
   337 => (x"48",x"d0",x"ff",x"b2"),
   338 => (x"73",x"78",x"e0",x"c0"),
   339 => (x"87",x"c2",x"02",x"9b"),
   340 => (x"48",x"75",x"7b",x"72"),
   341 => (x"4c",x"26",x"4d",x"26"),
   342 => (x"4f",x"26",x"4b",x"26"),
   343 => (x"0e",x"4f",x"26",x"1e"),
   344 => (x"0e",x"5c",x"5b",x"5e"),
   345 => (x"1e",x"76",x"86",x"f8"),
   346 => (x"fd",x"49",x"a6",x"c8"),
   347 => (x"86",x"c4",x"87",x"fd"),
   348 => (x"48",x"6e",x"4b",x"70"),
   349 => (x"c2",x"03",x"a8",x"c2"),
   350 => (x"4a",x"73",x"87",x"f0"),
   351 => (x"c1",x"9a",x"f0",x"c3"),
   352 => (x"c7",x"02",x"aa",x"d0"),
   353 => (x"aa",x"e0",x"c1",x"87"),
   354 => (x"87",x"de",x"c2",x"05"),
   355 => (x"99",x"c8",x"49",x"73"),
   356 => (x"ff",x"87",x"c3",x"02"),
   357 => (x"4c",x"73",x"87",x"c6"),
   358 => (x"ac",x"c2",x"9c",x"c3"),
   359 => (x"87",x"c2",x"c1",x"05"),
   360 => (x"c9",x"49",x"66",x"c4"),
   361 => (x"c4",x"1e",x"71",x"31"),
   362 => (x"92",x"d4",x"4a",x"66"),
   363 => (x"49",x"e1",x"ee",x"c2"),
   364 => (x"d0",x"fe",x"81",x"72"),
   365 => (x"49",x"d8",x"87",x"d1"),
   366 => (x"87",x"c3",x"d8",x"ff"),
   367 => (x"c2",x"1e",x"c0",x"c8"),
   368 => (x"fd",x"49",x"fe",x"dc"),
   369 => (x"ff",x"87",x"d7",x"ec"),
   370 => (x"e0",x"c0",x"48",x"d0"),
   371 => (x"fe",x"dc",x"c2",x"78"),
   372 => (x"4a",x"66",x"cc",x"1e"),
   373 => (x"ee",x"c2",x"92",x"d4"),
   374 => (x"81",x"72",x"49",x"e1"),
   375 => (x"87",x"d9",x"ce",x"fe"),
   376 => (x"ac",x"c1",x"86",x"cc"),
   377 => (x"87",x"c2",x"c1",x"05"),
   378 => (x"c9",x"49",x"66",x"c4"),
   379 => (x"c4",x"1e",x"71",x"31"),
   380 => (x"92",x"d4",x"4a",x"66"),
   381 => (x"49",x"e1",x"ee",x"c2"),
   382 => (x"cf",x"fe",x"81",x"72"),
   383 => (x"dc",x"c2",x"87",x"c9"),
   384 => (x"66",x"c8",x"1e",x"fe"),
   385 => (x"c2",x"92",x"d4",x"4a"),
   386 => (x"72",x"49",x"e1",x"ee"),
   387 => (x"da",x"cc",x"fe",x"81"),
   388 => (x"ff",x"49",x"d7",x"87"),
   389 => (x"c8",x"87",x"e8",x"d6"),
   390 => (x"dc",x"c2",x"1e",x"c0"),
   391 => (x"ea",x"fd",x"49",x"fe"),
   392 => (x"86",x"cc",x"87",x"d5"),
   393 => (x"c0",x"48",x"d0",x"ff"),
   394 => (x"8e",x"f8",x"78",x"e0"),
   395 => (x"0e",x"87",x"e7",x"fc"),
   396 => (x"5d",x"5c",x"5b",x"5e"),
   397 => (x"4d",x"71",x"1e",x"0e"),
   398 => (x"d4",x"4c",x"d4",x"ff"),
   399 => (x"c3",x"48",x"7e",x"66"),
   400 => (x"c5",x"06",x"a8",x"b7"),
   401 => (x"c1",x"48",x"c0",x"87"),
   402 => (x"49",x"75",x"87",x"e9"),
   403 => (x"87",x"ff",x"dc",x"fe"),
   404 => (x"66",x"c4",x"1e",x"75"),
   405 => (x"c2",x"93",x"d4",x"4b"),
   406 => (x"73",x"83",x"e1",x"ee"),
   407 => (x"d8",x"c6",x"fe",x"49"),
   408 => (x"6b",x"83",x"c8",x"87"),
   409 => (x"48",x"d0",x"ff",x"4b"),
   410 => (x"dd",x"78",x"e1",x"c8"),
   411 => (x"c3",x"48",x"73",x"7c"),
   412 => (x"7c",x"70",x"98",x"ff"),
   413 => (x"b7",x"c8",x"49",x"73"),
   414 => (x"c3",x"48",x"71",x"29"),
   415 => (x"7c",x"70",x"98",x"ff"),
   416 => (x"b7",x"d0",x"49",x"73"),
   417 => (x"c3",x"48",x"71",x"29"),
   418 => (x"7c",x"70",x"98",x"ff"),
   419 => (x"b7",x"d8",x"48",x"73"),
   420 => (x"c0",x"7c",x"70",x"28"),
   421 => (x"7c",x"7c",x"7c",x"7c"),
   422 => (x"7c",x"7c",x"7c",x"7c"),
   423 => (x"7c",x"7c",x"7c",x"7c"),
   424 => (x"c0",x"48",x"d0",x"ff"),
   425 => (x"66",x"c4",x"78",x"e0"),
   426 => (x"ff",x"49",x"dc",x"1e"),
   427 => (x"c8",x"87",x"f5",x"d4"),
   428 => (x"26",x"48",x"73",x"86"),
   429 => (x"1e",x"87",x"dd",x"fa"),
   430 => (x"4b",x"c0",x"1e",x"73"),
   431 => (x"f8",x"db",x"c2",x"1e"),
   432 => (x"ea",x"fd",x"49",x"bf"),
   433 => (x"c2",x"86",x"c4",x"87"),
   434 => (x"49",x"bf",x"fc",x"db"),
   435 => (x"87",x"e3",x"de",x"fe"),
   436 => (x"c4",x"05",x"98",x"70"),
   437 => (x"e5",x"db",x"c2",x"87"),
   438 => (x"c4",x"48",x"73",x"4b"),
   439 => (x"26",x"4d",x"26",x"87"),
   440 => (x"26",x"4b",x"26",x"4c"),
   441 => (x"4d",x"4f",x"52",x"4f"),
   442 => (x"61",x"6f",x"6c",x"20"),
   443 => (x"67",x"6e",x"69",x"64"),
   444 => (x"69",x"61",x"66",x"20"),
   445 => (x"00",x"64",x"65",x"6c"),
   446 => (x"00",x"00",x"27",x"00"),
   447 => (x"00",x"00",x"27",x"0c"),
   448 => (x"20",x"43",x"42",x"42"),
   449 => (x"20",x"20",x"20",x"20"),
   450 => (x"00",x"44",x"48",x"56"),
   451 => (x"20",x"43",x"42",x"42"),
   452 => (x"20",x"20",x"20",x"20"),
   453 => (x"00",x"4d",x"4f",x"52"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

