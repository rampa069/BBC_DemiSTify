
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c4",x"f6",x"c2",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"c4",x"f6",x"c2"),
    18 => (x"48",x"cc",x"e3",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"cc",x"e3",x"c2",x"87"),
    25 => (x"c8",x"e3",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e8",x"c1",x"87",x"f7"),
    29 => (x"e3",x"c2",x"87",x"c2"),
    30 => (x"e3",x"c2",x"4d",x"cc"),
    31 => (x"ad",x"74",x"4c",x"cc"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"73",x"1e",x"74",x"1e"),
    65 => (x"c1",x"1e",x"72",x"1e"),
    66 => (x"87",x"d0",x"04",x"8b"),
    67 => (x"02",x"11",x"48",x"12"),
    68 => (x"c3",x"4c",x"87",x"ca"),
    69 => (x"74",x"9c",x"98",x"df"),
    70 => (x"87",x"eb",x"02",x"88"),
    71 => (x"4b",x"26",x"4a",x"26"),
    72 => (x"4f",x"26",x"4c",x"26"),
    73 => (x"81",x"48",x"73",x"1e"),
    74 => (x"c5",x"02",x"a9",x"73"),
    75 => (x"05",x"53",x"12",x"87"),
    76 => (x"4f",x"26",x"87",x"f6"),
    77 => (x"71",x"1e",x"73",x"1e"),
    78 => (x"4b",x"66",x"c8",x"4a"),
    79 => (x"71",x"8b",x"c1",x"49"),
    80 => (x"87",x"cf",x"02",x"99"),
    81 => (x"d4",x"ff",x"48",x"12"),
    82 => (x"49",x"73",x"78",x"08"),
    83 => (x"99",x"71",x"8b",x"c1"),
    84 => (x"26",x"87",x"f1",x"05"),
    85 => (x"0e",x"4f",x"26",x"4b"),
    86 => (x"0e",x"5c",x"5b",x"5e"),
    87 => (x"d4",x"ff",x"4a",x"71"),
    88 => (x"4b",x"66",x"cc",x"4c"),
    89 => (x"71",x"8b",x"c1",x"49"),
    90 => (x"87",x"ce",x"02",x"99"),
    91 => (x"6c",x"7c",x"ff",x"c3"),
    92 => (x"c1",x"49",x"73",x"52"),
    93 => (x"05",x"99",x"71",x"8b"),
    94 => (x"4c",x"26",x"87",x"f2"),
    95 => (x"4f",x"26",x"4b",x"26"),
    96 => (x"ff",x"1e",x"73",x"1e"),
    97 => (x"ff",x"c3",x"4b",x"d4"),
    98 => (x"c3",x"4a",x"6b",x"7b"),
    99 => (x"49",x"6b",x"7b",x"ff"),
   100 => (x"b1",x"72",x"32",x"c8"),
   101 => (x"6b",x"7b",x"ff",x"c3"),
   102 => (x"71",x"31",x"c8",x"4a"),
   103 => (x"7b",x"ff",x"c3",x"b2"),
   104 => (x"32",x"c8",x"49",x"6b"),
   105 => (x"48",x"71",x"b1",x"72"),
   106 => (x"4f",x"26",x"4b",x"26"),
   107 => (x"5c",x"5b",x"5e",x"0e"),
   108 => (x"4d",x"71",x"0e",x"5d"),
   109 => (x"75",x"4c",x"d4",x"ff"),
   110 => (x"98",x"ff",x"c3",x"48"),
   111 => (x"e3",x"c2",x"7c",x"70"),
   112 => (x"c8",x"05",x"bf",x"cc"),
   113 => (x"48",x"66",x"d0",x"87"),
   114 => (x"a6",x"d4",x"30",x"c9"),
   115 => (x"49",x"66",x"d0",x"58"),
   116 => (x"48",x"71",x"29",x"d8"),
   117 => (x"70",x"98",x"ff",x"c3"),
   118 => (x"49",x"66",x"d0",x"7c"),
   119 => (x"48",x"71",x"29",x"d0"),
   120 => (x"70",x"98",x"ff",x"c3"),
   121 => (x"49",x"66",x"d0",x"7c"),
   122 => (x"48",x"71",x"29",x"c8"),
   123 => (x"70",x"98",x"ff",x"c3"),
   124 => (x"48",x"66",x"d0",x"7c"),
   125 => (x"70",x"98",x"ff",x"c3"),
   126 => (x"d0",x"49",x"75",x"7c"),
   127 => (x"c3",x"48",x"71",x"29"),
   128 => (x"7c",x"70",x"98",x"ff"),
   129 => (x"f0",x"c9",x"4b",x"6c"),
   130 => (x"ff",x"c3",x"4a",x"ff"),
   131 => (x"87",x"cf",x"05",x"ab"),
   132 => (x"6c",x"7c",x"71",x"49"),
   133 => (x"02",x"8a",x"c1",x"4b"),
   134 => (x"ab",x"71",x"87",x"c5"),
   135 => (x"73",x"87",x"f2",x"02"),
   136 => (x"26",x"4d",x"26",x"48"),
   137 => (x"26",x"4b",x"26",x"4c"),
   138 => (x"49",x"c0",x"1e",x"4f"),
   139 => (x"c3",x"48",x"d4",x"ff"),
   140 => (x"81",x"c1",x"78",x"ff"),
   141 => (x"a9",x"b7",x"c8",x"c3"),
   142 => (x"26",x"87",x"f1",x"04"),
   143 => (x"5b",x"5e",x"0e",x"4f"),
   144 => (x"c0",x"0e",x"5d",x"5c"),
   145 => (x"f7",x"c1",x"f0",x"ff"),
   146 => (x"c0",x"c0",x"c1",x"4d"),
   147 => (x"4b",x"c0",x"c0",x"c0"),
   148 => (x"c4",x"87",x"d6",x"ff"),
   149 => (x"c0",x"4c",x"df",x"f8"),
   150 => (x"fd",x"49",x"75",x"1e"),
   151 => (x"86",x"c4",x"87",x"ce"),
   152 => (x"c0",x"05",x"a8",x"c1"),
   153 => (x"d4",x"ff",x"87",x"e5"),
   154 => (x"78",x"ff",x"c3",x"48"),
   155 => (x"e1",x"c0",x"1e",x"73"),
   156 => (x"49",x"e9",x"c1",x"f0"),
   157 => (x"c4",x"87",x"f5",x"fc"),
   158 => (x"05",x"98",x"70",x"86"),
   159 => (x"d4",x"ff",x"87",x"ca"),
   160 => (x"78",x"ff",x"c3",x"48"),
   161 => (x"87",x"cb",x"48",x"c1"),
   162 => (x"c1",x"87",x"de",x"fe"),
   163 => (x"c6",x"ff",x"05",x"8c"),
   164 => (x"26",x"48",x"c0",x"87"),
   165 => (x"26",x"4c",x"26",x"4d"),
   166 => (x"0e",x"4f",x"26",x"4b"),
   167 => (x"0e",x"5c",x"5b",x"5e"),
   168 => (x"c1",x"f0",x"ff",x"c0"),
   169 => (x"d4",x"ff",x"4c",x"c1"),
   170 => (x"78",x"ff",x"c3",x"48"),
   171 => (x"f7",x"49",x"e0",x"cb"),
   172 => (x"4b",x"d3",x"87",x"f5"),
   173 => (x"49",x"74",x"1e",x"c0"),
   174 => (x"c4",x"87",x"f1",x"fb"),
   175 => (x"05",x"98",x"70",x"86"),
   176 => (x"d4",x"ff",x"87",x"ca"),
   177 => (x"78",x"ff",x"c3",x"48"),
   178 => (x"87",x"cb",x"48",x"c1"),
   179 => (x"c1",x"87",x"da",x"fd"),
   180 => (x"df",x"ff",x"05",x"8b"),
   181 => (x"26",x"48",x"c0",x"87"),
   182 => (x"26",x"4b",x"26",x"4c"),
   183 => (x"00",x"00",x"00",x"4f"),
   184 => (x"00",x"44",x"4d",x"43"),
   185 => (x"5c",x"5b",x"5e",x"0e"),
   186 => (x"ff",x"c3",x"0e",x"5d"),
   187 => (x"4b",x"d4",x"ff",x"4d"),
   188 => (x"c6",x"87",x"f6",x"fc"),
   189 => (x"e1",x"c0",x"1e",x"ea"),
   190 => (x"49",x"c8",x"c1",x"f0"),
   191 => (x"c4",x"87",x"ed",x"fa"),
   192 => (x"02",x"a8",x"c1",x"86"),
   193 => (x"d2",x"fe",x"87",x"c8"),
   194 => (x"c1",x"48",x"c0",x"87"),
   195 => (x"ef",x"f9",x"87",x"e8"),
   196 => (x"cf",x"49",x"70",x"87"),
   197 => (x"c6",x"99",x"ff",x"ff"),
   198 => (x"c8",x"02",x"a9",x"ea"),
   199 => (x"87",x"fb",x"fd",x"87"),
   200 => (x"d1",x"c1",x"48",x"c0"),
   201 => (x"c0",x"7b",x"75",x"87"),
   202 => (x"d0",x"fc",x"4c",x"f1"),
   203 => (x"02",x"98",x"70",x"87"),
   204 => (x"c0",x"87",x"ec",x"c0"),
   205 => (x"f0",x"ff",x"c0",x"1e"),
   206 => (x"f9",x"49",x"fa",x"c1"),
   207 => (x"86",x"c4",x"87",x"ee"),
   208 => (x"da",x"05",x"98",x"70"),
   209 => (x"6b",x"7b",x"75",x"87"),
   210 => (x"75",x"7b",x"75",x"49"),
   211 => (x"75",x"7b",x"75",x"7b"),
   212 => (x"99",x"c0",x"c1",x"7b"),
   213 => (x"c1",x"87",x"c4",x"02"),
   214 => (x"c0",x"87",x"db",x"48"),
   215 => (x"c2",x"87",x"d7",x"48"),
   216 => (x"87",x"ca",x"05",x"ac"),
   217 => (x"f4",x"49",x"c0",x"ce"),
   218 => (x"48",x"c0",x"87",x"fd"),
   219 => (x"8c",x"c1",x"87",x"c8"),
   220 => (x"87",x"f6",x"fe",x"05"),
   221 => (x"4d",x"26",x"48",x"c0"),
   222 => (x"4b",x"26",x"4c",x"26"),
   223 => (x"00",x"00",x"4f",x"26"),
   224 => (x"43",x"48",x"44",x"53"),
   225 => (x"69",x"61",x"66",x"20"),
   226 => (x"00",x"0a",x"21",x"6c"),
   227 => (x"5c",x"5b",x"5e",x"0e"),
   228 => (x"d0",x"ff",x"0e",x"5d"),
   229 => (x"d0",x"e5",x"c0",x"4d"),
   230 => (x"c2",x"4c",x"c0",x"c1"),
   231 => (x"c1",x"48",x"cc",x"e3"),
   232 => (x"49",x"d8",x"d0",x"78"),
   233 => (x"c7",x"87",x"c0",x"f4"),
   234 => (x"f9",x"7d",x"c2",x"4b"),
   235 => (x"7d",x"c3",x"87",x"fb"),
   236 => (x"49",x"74",x"1e",x"c0"),
   237 => (x"c4",x"87",x"f5",x"f7"),
   238 => (x"05",x"a8",x"c1",x"86"),
   239 => (x"c2",x"4b",x"87",x"c1"),
   240 => (x"87",x"cb",x"05",x"ab"),
   241 => (x"f3",x"49",x"d0",x"d0"),
   242 => (x"48",x"c0",x"87",x"dd"),
   243 => (x"c1",x"87",x"f6",x"c0"),
   244 => (x"d4",x"ff",x"05",x"8b"),
   245 => (x"87",x"cc",x"fc",x"87"),
   246 => (x"58",x"d0",x"e3",x"c2"),
   247 => (x"cd",x"05",x"98",x"70"),
   248 => (x"c0",x"1e",x"c1",x"87"),
   249 => (x"d0",x"c1",x"f0",x"ff"),
   250 => (x"87",x"c0",x"f7",x"49"),
   251 => (x"d4",x"ff",x"86",x"c4"),
   252 => (x"78",x"ff",x"c3",x"48"),
   253 => (x"c2",x"87",x"cc",x"c5"),
   254 => (x"c2",x"58",x"d4",x"e3"),
   255 => (x"48",x"d4",x"ff",x"7d"),
   256 => (x"c1",x"78",x"ff",x"c3"),
   257 => (x"26",x"4d",x"26",x"48"),
   258 => (x"26",x"4b",x"26",x"4c"),
   259 => (x"00",x"00",x"00",x"4f"),
   260 => (x"52",x"52",x"45",x"49"),
   261 => (x"00",x"00",x"00",x"00"),
   262 => (x"00",x"49",x"50",x"53"),
   263 => (x"5c",x"5b",x"5e",x"0e"),
   264 => (x"4d",x"71",x"0e",x"5d"),
   265 => (x"ff",x"4c",x"ff",x"c3"),
   266 => (x"7b",x"74",x"4b",x"d4"),
   267 => (x"c4",x"48",x"d0",x"ff"),
   268 => (x"7b",x"74",x"78",x"c3"),
   269 => (x"ff",x"c0",x"1e",x"75"),
   270 => (x"49",x"d8",x"c1",x"f0"),
   271 => (x"c4",x"87",x"ed",x"f5"),
   272 => (x"02",x"98",x"70",x"86"),
   273 => (x"c8",x"d2",x"87",x"cb"),
   274 => (x"87",x"db",x"f1",x"49"),
   275 => (x"ee",x"c0",x"48",x"c1"),
   276 => (x"c3",x"7b",x"74",x"87"),
   277 => (x"c0",x"c8",x"7b",x"fe"),
   278 => (x"49",x"66",x"d4",x"1e"),
   279 => (x"c4",x"87",x"d5",x"f3"),
   280 => (x"74",x"7b",x"74",x"86"),
   281 => (x"d8",x"7b",x"74",x"7b"),
   282 => (x"74",x"4a",x"e0",x"da"),
   283 => (x"c5",x"05",x"6b",x"7b"),
   284 => (x"05",x"8a",x"c1",x"87"),
   285 => (x"7b",x"74",x"87",x"f5"),
   286 => (x"c2",x"48",x"d0",x"ff"),
   287 => (x"26",x"48",x"c0",x"78"),
   288 => (x"26",x"4c",x"26",x"4d"),
   289 => (x"00",x"4f",x"26",x"4b"),
   290 => (x"74",x"69",x"72",x"57"),
   291 => (x"61",x"66",x"20",x"65"),
   292 => (x"64",x"65",x"6c",x"69"),
   293 => (x"5e",x"0e",x"00",x"0a"),
   294 => (x"0e",x"5d",x"5c",x"5b"),
   295 => (x"4b",x"71",x"86",x"fc"),
   296 => (x"c0",x"4c",x"d4",x"ff"),
   297 => (x"cd",x"ee",x"c5",x"7e"),
   298 => (x"ff",x"c3",x"4a",x"df"),
   299 => (x"c3",x"48",x"6c",x"7c"),
   300 => (x"c0",x"05",x"a8",x"fe"),
   301 => (x"4d",x"74",x"87",x"f8"),
   302 => (x"cc",x"02",x"9b",x"73"),
   303 => (x"1e",x"66",x"d4",x"87"),
   304 => (x"d2",x"f2",x"49",x"73"),
   305 => (x"d4",x"86",x"c4",x"87"),
   306 => (x"48",x"d0",x"ff",x"87"),
   307 => (x"d4",x"78",x"d1",x"c4"),
   308 => (x"ff",x"c3",x"4a",x"66"),
   309 => (x"05",x"8a",x"c1",x"7d"),
   310 => (x"a6",x"d8",x"87",x"f8"),
   311 => (x"7c",x"ff",x"c3",x"5a"),
   312 => (x"05",x"9b",x"73",x"7c"),
   313 => (x"d0",x"ff",x"87",x"c5"),
   314 => (x"c1",x"78",x"d0",x"48"),
   315 => (x"8a",x"c1",x"7e",x"4a"),
   316 => (x"87",x"f6",x"fe",x"05"),
   317 => (x"8e",x"fc",x"48",x"6e"),
   318 => (x"4c",x"26",x"4d",x"26"),
   319 => (x"4f",x"26",x"4b",x"26"),
   320 => (x"71",x"1e",x"73",x"1e"),
   321 => (x"ff",x"4b",x"c0",x"4a"),
   322 => (x"ff",x"c3",x"48",x"d4"),
   323 => (x"48",x"d0",x"ff",x"78"),
   324 => (x"ff",x"78",x"c3",x"c4"),
   325 => (x"ff",x"c3",x"48",x"d4"),
   326 => (x"c0",x"1e",x"72",x"78"),
   327 => (x"d1",x"c1",x"f0",x"ff"),
   328 => (x"87",x"c8",x"f2",x"49"),
   329 => (x"98",x"70",x"86",x"c4"),
   330 => (x"c8",x"87",x"d2",x"05"),
   331 => (x"66",x"cc",x"1e",x"c0"),
   332 => (x"87",x"e2",x"fd",x"49"),
   333 => (x"4b",x"70",x"86",x"c4"),
   334 => (x"c2",x"48",x"d0",x"ff"),
   335 => (x"26",x"48",x"73",x"78"),
   336 => (x"0e",x"4f",x"26",x"4b"),
   337 => (x"5d",x"5c",x"5b",x"5e"),
   338 => (x"c0",x"1e",x"c0",x"0e"),
   339 => (x"c9",x"c1",x"f0",x"ff"),
   340 => (x"87",x"d8",x"f1",x"49"),
   341 => (x"e3",x"c2",x"1e",x"d2"),
   342 => (x"f9",x"fc",x"49",x"d4"),
   343 => (x"c0",x"86",x"c8",x"87"),
   344 => (x"d2",x"84",x"c1",x"4c"),
   345 => (x"f8",x"04",x"ac",x"b7"),
   346 => (x"d4",x"e3",x"c2",x"87"),
   347 => (x"c3",x"49",x"bf",x"97"),
   348 => (x"c0",x"c1",x"99",x"c0"),
   349 => (x"e7",x"c0",x"05",x"a9"),
   350 => (x"db",x"e3",x"c2",x"87"),
   351 => (x"d0",x"49",x"bf",x"97"),
   352 => (x"dc",x"e3",x"c2",x"31"),
   353 => (x"c8",x"4a",x"bf",x"97"),
   354 => (x"c2",x"b1",x"72",x"32"),
   355 => (x"bf",x"97",x"dd",x"e3"),
   356 => (x"4c",x"71",x"b1",x"4a"),
   357 => (x"ff",x"ff",x"ff",x"cf"),
   358 => (x"ca",x"84",x"c1",x"9c"),
   359 => (x"87",x"e7",x"c1",x"34"),
   360 => (x"97",x"dd",x"e3",x"c2"),
   361 => (x"31",x"c1",x"49",x"bf"),
   362 => (x"e3",x"c2",x"99",x"c6"),
   363 => (x"4a",x"bf",x"97",x"de"),
   364 => (x"72",x"2a",x"b7",x"c7"),
   365 => (x"d9",x"e3",x"c2",x"b1"),
   366 => (x"4d",x"4a",x"bf",x"97"),
   367 => (x"e3",x"c2",x"9d",x"cf"),
   368 => (x"4a",x"bf",x"97",x"da"),
   369 => (x"32",x"ca",x"9a",x"c3"),
   370 => (x"97",x"db",x"e3",x"c2"),
   371 => (x"33",x"c2",x"4b",x"bf"),
   372 => (x"e3",x"c2",x"b2",x"73"),
   373 => (x"4b",x"bf",x"97",x"dc"),
   374 => (x"c6",x"9b",x"c0",x"c3"),
   375 => (x"b2",x"73",x"2b",x"b7"),
   376 => (x"48",x"c1",x"81",x"c2"),
   377 => (x"49",x"70",x"30",x"71"),
   378 => (x"30",x"75",x"48",x"c1"),
   379 => (x"4c",x"72",x"4d",x"70"),
   380 => (x"94",x"71",x"84",x"c1"),
   381 => (x"ad",x"b7",x"c0",x"c8"),
   382 => (x"c1",x"87",x"cc",x"06"),
   383 => (x"c8",x"2d",x"b7",x"34"),
   384 => (x"01",x"ad",x"b7",x"c0"),
   385 => (x"74",x"87",x"f4",x"ff"),
   386 => (x"26",x"4d",x"26",x"48"),
   387 => (x"26",x"4b",x"26",x"4c"),
   388 => (x"5b",x"5e",x"0e",x"4f"),
   389 => (x"f8",x"0e",x"5d",x"5c"),
   390 => (x"fc",x"eb",x"c2",x"86"),
   391 => (x"c2",x"78",x"c0",x"48"),
   392 => (x"c0",x"1e",x"f4",x"e3"),
   393 => (x"87",x"d8",x"fb",x"49"),
   394 => (x"98",x"70",x"86",x"c4"),
   395 => (x"c0",x"87",x"c5",x"05"),
   396 => (x"87",x"c0",x"c9",x"48"),
   397 => (x"7e",x"c1",x"4d",x"c0"),
   398 => (x"bf",x"d8",x"f7",x"c0"),
   399 => (x"ea",x"e4",x"c2",x"49"),
   400 => (x"4b",x"c8",x"71",x"4a"),
   401 => (x"70",x"87",x"df",x"ea"),
   402 => (x"87",x"c2",x"05",x"98"),
   403 => (x"f7",x"c0",x"7e",x"c0"),
   404 => (x"c2",x"49",x"bf",x"d4"),
   405 => (x"71",x"4a",x"c6",x"e5"),
   406 => (x"c9",x"ea",x"4b",x"c8"),
   407 => (x"05",x"98",x"70",x"87"),
   408 => (x"7e",x"c0",x"87",x"c2"),
   409 => (x"fd",x"c0",x"02",x"6e"),
   410 => (x"fa",x"ea",x"c2",x"87"),
   411 => (x"eb",x"c2",x"4d",x"bf"),
   412 => (x"7e",x"bf",x"9f",x"f2"),
   413 => (x"ea",x"d6",x"c5",x"48"),
   414 => (x"87",x"c7",x"05",x"a8"),
   415 => (x"bf",x"fa",x"ea",x"c2"),
   416 => (x"6e",x"87",x"ce",x"4d"),
   417 => (x"d5",x"e9",x"ca",x"48"),
   418 => (x"87",x"c5",x"02",x"a8"),
   419 => (x"e3",x"c7",x"48",x"c0"),
   420 => (x"f4",x"e3",x"c2",x"87"),
   421 => (x"f9",x"49",x"75",x"1e"),
   422 => (x"86",x"c4",x"87",x"e6"),
   423 => (x"c5",x"05",x"98",x"70"),
   424 => (x"c7",x"48",x"c0",x"87"),
   425 => (x"f7",x"c0",x"87",x"ce"),
   426 => (x"c2",x"49",x"bf",x"d4"),
   427 => (x"71",x"4a",x"c6",x"e5"),
   428 => (x"f1",x"e8",x"4b",x"c8"),
   429 => (x"05",x"98",x"70",x"87"),
   430 => (x"eb",x"c2",x"87",x"c8"),
   431 => (x"78",x"c1",x"48",x"fc"),
   432 => (x"f7",x"c0",x"87",x"da"),
   433 => (x"c2",x"49",x"bf",x"d8"),
   434 => (x"71",x"4a",x"ea",x"e4"),
   435 => (x"d5",x"e8",x"4b",x"c8"),
   436 => (x"02",x"98",x"70",x"87"),
   437 => (x"c0",x"87",x"c5",x"c0"),
   438 => (x"87",x"d8",x"c6",x"48"),
   439 => (x"97",x"f2",x"eb",x"c2"),
   440 => (x"d5",x"c1",x"49",x"bf"),
   441 => (x"cd",x"c0",x"05",x"a9"),
   442 => (x"f3",x"eb",x"c2",x"87"),
   443 => (x"c2",x"49",x"bf",x"97"),
   444 => (x"c0",x"02",x"a9",x"ea"),
   445 => (x"48",x"c0",x"87",x"c5"),
   446 => (x"c2",x"87",x"f9",x"c5"),
   447 => (x"bf",x"97",x"f4",x"e3"),
   448 => (x"e9",x"c3",x"48",x"7e"),
   449 => (x"ce",x"c0",x"02",x"a8"),
   450 => (x"c3",x"48",x"6e",x"87"),
   451 => (x"c0",x"02",x"a8",x"eb"),
   452 => (x"48",x"c0",x"87",x"c5"),
   453 => (x"c2",x"87",x"dd",x"c5"),
   454 => (x"bf",x"97",x"ff",x"e3"),
   455 => (x"c0",x"05",x"99",x"49"),
   456 => (x"e4",x"c2",x"87",x"cc"),
   457 => (x"49",x"bf",x"97",x"c0"),
   458 => (x"c0",x"02",x"a9",x"c2"),
   459 => (x"48",x"c0",x"87",x"c5"),
   460 => (x"c2",x"87",x"c1",x"c5"),
   461 => (x"bf",x"97",x"c1",x"e4"),
   462 => (x"f8",x"eb",x"c2",x"48"),
   463 => (x"48",x"4c",x"70",x"58"),
   464 => (x"eb",x"c2",x"88",x"c1"),
   465 => (x"e4",x"c2",x"58",x"fc"),
   466 => (x"49",x"bf",x"97",x"c2"),
   467 => (x"e4",x"c2",x"81",x"75"),
   468 => (x"4a",x"bf",x"97",x"c3"),
   469 => (x"a1",x"72",x"32",x"c8"),
   470 => (x"cc",x"f0",x"c2",x"7e"),
   471 => (x"c2",x"78",x"6e",x"48"),
   472 => (x"bf",x"97",x"c4",x"e4"),
   473 => (x"58",x"a6",x"c8",x"48"),
   474 => (x"bf",x"fc",x"eb",x"c2"),
   475 => (x"87",x"cf",x"c2",x"02"),
   476 => (x"bf",x"d4",x"f7",x"c0"),
   477 => (x"c6",x"e5",x"c2",x"49"),
   478 => (x"4b",x"c8",x"71",x"4a"),
   479 => (x"70",x"87",x"e7",x"e5"),
   480 => (x"c5",x"c0",x"02",x"98"),
   481 => (x"c3",x"48",x"c0",x"87"),
   482 => (x"eb",x"c2",x"87",x"ea"),
   483 => (x"c2",x"4c",x"bf",x"f4"),
   484 => (x"c2",x"5c",x"e0",x"f0"),
   485 => (x"bf",x"97",x"d9",x"e4"),
   486 => (x"c2",x"31",x"c8",x"49"),
   487 => (x"bf",x"97",x"d8",x"e4"),
   488 => (x"c2",x"49",x"a1",x"4a"),
   489 => (x"bf",x"97",x"da",x"e4"),
   490 => (x"72",x"32",x"d0",x"4a"),
   491 => (x"e4",x"c2",x"49",x"a1"),
   492 => (x"4a",x"bf",x"97",x"db"),
   493 => (x"a1",x"72",x"32",x"d8"),
   494 => (x"91",x"66",x"c4",x"49"),
   495 => (x"bf",x"cc",x"f0",x"c2"),
   496 => (x"d4",x"f0",x"c2",x"81"),
   497 => (x"e1",x"e4",x"c2",x"59"),
   498 => (x"c8",x"4a",x"bf",x"97"),
   499 => (x"e0",x"e4",x"c2",x"32"),
   500 => (x"a2",x"4b",x"bf",x"97"),
   501 => (x"e2",x"e4",x"c2",x"4a"),
   502 => (x"d0",x"4b",x"bf",x"97"),
   503 => (x"4a",x"a2",x"73",x"33"),
   504 => (x"97",x"e3",x"e4",x"c2"),
   505 => (x"9b",x"cf",x"4b",x"bf"),
   506 => (x"a2",x"73",x"33",x"d8"),
   507 => (x"d8",x"f0",x"c2",x"4a"),
   508 => (x"74",x"8a",x"c2",x"5a"),
   509 => (x"d8",x"f0",x"c2",x"92"),
   510 => (x"78",x"a1",x"72",x"48"),
   511 => (x"c2",x"87",x"c1",x"c1"),
   512 => (x"bf",x"97",x"c6",x"e4"),
   513 => (x"c2",x"31",x"c8",x"49"),
   514 => (x"bf",x"97",x"c5",x"e4"),
   515 => (x"c5",x"49",x"a1",x"4a"),
   516 => (x"81",x"ff",x"c7",x"31"),
   517 => (x"f0",x"c2",x"29",x"c9"),
   518 => (x"e4",x"c2",x"59",x"e0"),
   519 => (x"4a",x"bf",x"97",x"cb"),
   520 => (x"e4",x"c2",x"32",x"c8"),
   521 => (x"4b",x"bf",x"97",x"ca"),
   522 => (x"66",x"c4",x"4a",x"a2"),
   523 => (x"c2",x"82",x"6e",x"92"),
   524 => (x"c2",x"5a",x"dc",x"f0"),
   525 => (x"c0",x"48",x"d4",x"f0"),
   526 => (x"d0",x"f0",x"c2",x"78"),
   527 => (x"78",x"a1",x"72",x"48"),
   528 => (x"48",x"e0",x"f0",x"c2"),
   529 => (x"bf",x"d4",x"f0",x"c2"),
   530 => (x"e4",x"f0",x"c2",x"78"),
   531 => (x"d8",x"f0",x"c2",x"48"),
   532 => (x"eb",x"c2",x"78",x"bf"),
   533 => (x"c0",x"02",x"bf",x"fc"),
   534 => (x"48",x"74",x"87",x"c9"),
   535 => (x"7e",x"70",x"30",x"c4"),
   536 => (x"c2",x"87",x"c9",x"c0"),
   537 => (x"48",x"bf",x"dc",x"f0"),
   538 => (x"7e",x"70",x"30",x"c4"),
   539 => (x"48",x"c0",x"ec",x"c2"),
   540 => (x"48",x"c1",x"78",x"6e"),
   541 => (x"4d",x"26",x"8e",x"f8"),
   542 => (x"4b",x"26",x"4c",x"26"),
   543 => (x"5e",x"0e",x"4f",x"26"),
   544 => (x"0e",x"5d",x"5c",x"5b"),
   545 => (x"eb",x"c2",x"4a",x"71"),
   546 => (x"cb",x"02",x"bf",x"fc"),
   547 => (x"c7",x"4b",x"72",x"87"),
   548 => (x"c1",x"4d",x"72",x"2b"),
   549 => (x"87",x"c9",x"9d",x"ff"),
   550 => (x"2b",x"c8",x"4b",x"72"),
   551 => (x"ff",x"c3",x"4d",x"72"),
   552 => (x"cc",x"f0",x"c2",x"9d"),
   553 => (x"f7",x"c0",x"83",x"bf"),
   554 => (x"02",x"ab",x"bf",x"d0"),
   555 => (x"f7",x"c0",x"87",x"d9"),
   556 => (x"e3",x"c2",x"5b",x"d4"),
   557 => (x"49",x"73",x"1e",x"f4"),
   558 => (x"c4",x"87",x"c5",x"f1"),
   559 => (x"05",x"98",x"70",x"86"),
   560 => (x"48",x"c0",x"87",x"c5"),
   561 => (x"c2",x"87",x"e6",x"c0"),
   562 => (x"02",x"bf",x"fc",x"eb"),
   563 => (x"49",x"75",x"87",x"d2"),
   564 => (x"e3",x"c2",x"91",x"c4"),
   565 => (x"4c",x"69",x"81",x"f4"),
   566 => (x"ff",x"ff",x"ff",x"cf"),
   567 => (x"87",x"cb",x"9c",x"ff"),
   568 => (x"91",x"c2",x"49",x"75"),
   569 => (x"81",x"f4",x"e3",x"c2"),
   570 => (x"74",x"4c",x"69",x"9f"),
   571 => (x"26",x"4d",x"26",x"48"),
   572 => (x"26",x"4b",x"26",x"4c"),
   573 => (x"5b",x"5e",x"0e",x"4f"),
   574 => (x"f4",x"0e",x"5d",x"5c"),
   575 => (x"59",x"a6",x"cc",x"86"),
   576 => (x"c5",x"05",x"66",x"c8"),
   577 => (x"c3",x"48",x"c0",x"87"),
   578 => (x"66",x"c8",x"87",x"c7"),
   579 => (x"70",x"80",x"c8",x"48"),
   580 => (x"78",x"c0",x"48",x"7e"),
   581 => (x"c7",x"02",x"66",x"dc"),
   582 => (x"97",x"66",x"dc",x"87"),
   583 => (x"87",x"c5",x"05",x"bf"),
   584 => (x"ec",x"c2",x"48",x"c0"),
   585 => (x"c1",x"1e",x"c0",x"87"),
   586 => (x"e9",x"ca",x"49",x"49"),
   587 => (x"70",x"86",x"c4",x"87"),
   588 => (x"c0",x"02",x"9c",x"4c"),
   589 => (x"ec",x"c2",x"87",x"fc"),
   590 => (x"66",x"dc",x"4a",x"c4"),
   591 => (x"ca",x"de",x"ff",x"49"),
   592 => (x"02",x"98",x"70",x"87"),
   593 => (x"74",x"87",x"eb",x"c0"),
   594 => (x"49",x"66",x"dc",x"4a"),
   595 => (x"de",x"ff",x"4b",x"cb"),
   596 => (x"98",x"70",x"87",x"ee"),
   597 => (x"c0",x"87",x"db",x"02"),
   598 => (x"02",x"9c",x"74",x"1e"),
   599 => (x"4d",x"c0",x"87",x"c4"),
   600 => (x"4d",x"c1",x"87",x"c2"),
   601 => (x"ed",x"c9",x"49",x"75"),
   602 => (x"70",x"86",x"c4",x"87"),
   603 => (x"ff",x"05",x"9c",x"4c"),
   604 => (x"9c",x"74",x"87",x"c4"),
   605 => (x"87",x"d7",x"c1",x"02"),
   606 => (x"6e",x"49",x"a4",x"dc"),
   607 => (x"da",x"78",x"69",x"48"),
   608 => (x"66",x"c8",x"49",x"a4"),
   609 => (x"c8",x"80",x"c4",x"48"),
   610 => (x"69",x"9f",x"58",x"a6"),
   611 => (x"08",x"66",x"c4",x"48"),
   612 => (x"fc",x"eb",x"c2",x"78"),
   613 => (x"87",x"d2",x"02",x"bf"),
   614 => (x"9f",x"49",x"a4",x"d4"),
   615 => (x"ff",x"c0",x"49",x"69"),
   616 => (x"48",x"71",x"99",x"ff"),
   617 => (x"7e",x"70",x"30",x"d0"),
   618 => (x"7e",x"c0",x"87",x"c2"),
   619 => (x"66",x"c4",x"48",x"6e"),
   620 => (x"66",x"c4",x"80",x"bf"),
   621 => (x"66",x"c8",x"78",x"08"),
   622 => (x"c8",x"78",x"c0",x"48"),
   623 => (x"81",x"cc",x"49",x"66"),
   624 => (x"79",x"bf",x"66",x"c4"),
   625 => (x"d0",x"49",x"66",x"c8"),
   626 => (x"c1",x"79",x"c0",x"81"),
   627 => (x"c0",x"87",x"c2",x"48"),
   628 => (x"26",x"8e",x"f4",x"48"),
   629 => (x"26",x"4c",x"26",x"4d"),
   630 => (x"0e",x"4f",x"26",x"4b"),
   631 => (x"5d",x"5c",x"5b",x"5e"),
   632 => (x"d0",x"4c",x"71",x"0e"),
   633 => (x"9c",x"74",x"4d",x"66"),
   634 => (x"87",x"c2",x"c1",x"02"),
   635 => (x"69",x"49",x"a4",x"c8"),
   636 => (x"87",x"fa",x"c0",x"02"),
   637 => (x"75",x"85",x"49",x"6c"),
   638 => (x"f8",x"eb",x"c2",x"b9"),
   639 => (x"ba",x"ff",x"4a",x"bf"),
   640 => (x"99",x"71",x"99",x"72"),
   641 => (x"87",x"e4",x"c0",x"02"),
   642 => (x"6b",x"4b",x"a4",x"c4"),
   643 => (x"87",x"ee",x"f9",x"49"),
   644 => (x"eb",x"c2",x"7b",x"70"),
   645 => (x"6c",x"49",x"bf",x"f4"),
   646 => (x"75",x"7c",x"71",x"81"),
   647 => (x"f8",x"eb",x"c2",x"b9"),
   648 => (x"ba",x"ff",x"4a",x"bf"),
   649 => (x"99",x"71",x"99",x"72"),
   650 => (x"87",x"dc",x"ff",x"05"),
   651 => (x"4d",x"26",x"7c",x"75"),
   652 => (x"4b",x"26",x"4c",x"26"),
   653 => (x"73",x"1e",x"4f",x"26"),
   654 => (x"9b",x"4b",x"71",x"1e"),
   655 => (x"c8",x"87",x"c7",x"02"),
   656 => (x"05",x"69",x"49",x"a3"),
   657 => (x"48",x"c0",x"87",x"c5"),
   658 => (x"c2",x"87",x"f6",x"c0"),
   659 => (x"49",x"bf",x"d0",x"f0"),
   660 => (x"6a",x"4a",x"a3",x"c4"),
   661 => (x"c2",x"8a",x"c2",x"4a"),
   662 => (x"92",x"bf",x"f4",x"eb"),
   663 => (x"c2",x"49",x"a1",x"72"),
   664 => (x"4a",x"bf",x"f8",x"eb"),
   665 => (x"a1",x"72",x"9a",x"6b"),
   666 => (x"d4",x"f7",x"c0",x"49"),
   667 => (x"1e",x"66",x"c8",x"59"),
   668 => (x"87",x"cc",x"ea",x"71"),
   669 => (x"98",x"70",x"86",x"c4"),
   670 => (x"c0",x"87",x"c4",x"05"),
   671 => (x"c1",x"87",x"c2",x"48"),
   672 => (x"26",x"4b",x"26",x"48"),
   673 => (x"1e",x"73",x"1e",x"4f"),
   674 => (x"02",x"9b",x"4b",x"71"),
   675 => (x"a3",x"c8",x"87",x"c7"),
   676 => (x"c5",x"05",x"69",x"49"),
   677 => (x"c0",x"48",x"c0",x"87"),
   678 => (x"f0",x"c2",x"87",x"f6"),
   679 => (x"c4",x"49",x"bf",x"d0"),
   680 => (x"4a",x"6a",x"4a",x"a3"),
   681 => (x"eb",x"c2",x"8a",x"c2"),
   682 => (x"72",x"92",x"bf",x"f4"),
   683 => (x"eb",x"c2",x"49",x"a1"),
   684 => (x"6b",x"4a",x"bf",x"f8"),
   685 => (x"49",x"a1",x"72",x"9a"),
   686 => (x"59",x"d4",x"f7",x"c0"),
   687 => (x"71",x"1e",x"66",x"c8"),
   688 => (x"c4",x"87",x"d9",x"e5"),
   689 => (x"05",x"98",x"70",x"86"),
   690 => (x"48",x"c0",x"87",x"c4"),
   691 => (x"48",x"c1",x"87",x"c2"),
   692 => (x"4f",x"26",x"4b",x"26"),
   693 => (x"5c",x"5b",x"5e",x"0e"),
   694 => (x"86",x"fc",x"0e",x"5d"),
   695 => (x"66",x"d4",x"4b",x"71"),
   696 => (x"02",x"9b",x"73",x"4d"),
   697 => (x"c8",x"87",x"cc",x"c1"),
   698 => (x"02",x"69",x"49",x"a3"),
   699 => (x"d0",x"87",x"c4",x"c1"),
   700 => (x"eb",x"c2",x"4c",x"a3"),
   701 => (x"ff",x"49",x"bf",x"f8"),
   702 => (x"99",x"4a",x"6c",x"b9"),
   703 => (x"a9",x"66",x"d4",x"7e"),
   704 => (x"c0",x"87",x"cd",x"06"),
   705 => (x"a3",x"cc",x"7c",x"7b"),
   706 => (x"49",x"a3",x"c4",x"4a"),
   707 => (x"87",x"ca",x"79",x"6a"),
   708 => (x"c0",x"f8",x"49",x"72"),
   709 => (x"4d",x"66",x"d4",x"99"),
   710 => (x"49",x"75",x"8d",x"71"),
   711 => (x"1e",x"71",x"29",x"c9"),
   712 => (x"f6",x"fa",x"49",x"73"),
   713 => (x"f4",x"e3",x"c2",x"87"),
   714 => (x"fc",x"49",x"73",x"1e"),
   715 => (x"86",x"c8",x"87",x"c8"),
   716 => (x"fc",x"7c",x"66",x"d4"),
   717 => (x"26",x"4d",x"26",x"8e"),
   718 => (x"26",x"4b",x"26",x"4c"),
   719 => (x"1e",x"73",x"1e",x"4f"),
   720 => (x"02",x"9b",x"4b",x"71"),
   721 => (x"c2",x"87",x"e4",x"c0"),
   722 => (x"73",x"5b",x"e4",x"f0"),
   723 => (x"c2",x"8a",x"c2",x"4a"),
   724 => (x"49",x"bf",x"f4",x"eb"),
   725 => (x"d0",x"f0",x"c2",x"92"),
   726 => (x"80",x"72",x"48",x"bf"),
   727 => (x"58",x"e8",x"f0",x"c2"),
   728 => (x"30",x"c4",x"48",x"71"),
   729 => (x"58",x"c4",x"ec",x"c2"),
   730 => (x"c2",x"87",x"ed",x"c0"),
   731 => (x"c2",x"48",x"e0",x"f0"),
   732 => (x"78",x"bf",x"d4",x"f0"),
   733 => (x"48",x"e4",x"f0",x"c2"),
   734 => (x"bf",x"d8",x"f0",x"c2"),
   735 => (x"fc",x"eb",x"c2",x"78"),
   736 => (x"87",x"c9",x"02",x"bf"),
   737 => (x"bf",x"f4",x"eb",x"c2"),
   738 => (x"c7",x"31",x"c4",x"49"),
   739 => (x"dc",x"f0",x"c2",x"87"),
   740 => (x"31",x"c4",x"49",x"bf"),
   741 => (x"59",x"c4",x"ec",x"c2"),
   742 => (x"4f",x"26",x"4b",x"26"),
   743 => (x"5c",x"5b",x"5e",x"0e"),
   744 => (x"c0",x"4a",x"71",x"0e"),
   745 => (x"02",x"9a",x"72",x"4b"),
   746 => (x"da",x"87",x"e0",x"c0"),
   747 => (x"69",x"9f",x"49",x"a2"),
   748 => (x"fc",x"eb",x"c2",x"4b"),
   749 => (x"87",x"cf",x"02",x"bf"),
   750 => (x"9f",x"49",x"a2",x"d4"),
   751 => (x"c0",x"4c",x"49",x"69"),
   752 => (x"d0",x"9c",x"ff",x"ff"),
   753 => (x"c0",x"87",x"c2",x"34"),
   754 => (x"73",x"b3",x"74",x"4c"),
   755 => (x"87",x"ed",x"fd",x"49"),
   756 => (x"4b",x"26",x"4c",x"26"),
   757 => (x"5e",x"0e",x"4f",x"26"),
   758 => (x"0e",x"5d",x"5c",x"5b"),
   759 => (x"a6",x"c8",x"86",x"f0"),
   760 => (x"ff",x"ff",x"cf",x"59"),
   761 => (x"c0",x"4c",x"f8",x"ff"),
   762 => (x"02",x"66",x"c4",x"7e"),
   763 => (x"e3",x"c2",x"87",x"d8"),
   764 => (x"78",x"c0",x"48",x"f0"),
   765 => (x"48",x"e8",x"e3",x"c2"),
   766 => (x"bf",x"e4",x"f0",x"c2"),
   767 => (x"ec",x"e3",x"c2",x"78"),
   768 => (x"e0",x"f0",x"c2",x"48"),
   769 => (x"ec",x"c2",x"78",x"bf"),
   770 => (x"50",x"c0",x"48",x"d1"),
   771 => (x"bf",x"c0",x"ec",x"c2"),
   772 => (x"f0",x"e3",x"c2",x"49"),
   773 => (x"aa",x"71",x"4a",x"bf"),
   774 => (x"87",x"cb",x"c4",x"03"),
   775 => (x"99",x"cf",x"49",x"72"),
   776 => (x"87",x"e9",x"c0",x"05"),
   777 => (x"48",x"d0",x"f7",x"c0"),
   778 => (x"bf",x"e8",x"e3",x"c2"),
   779 => (x"f4",x"e3",x"c2",x"78"),
   780 => (x"e8",x"e3",x"c2",x"1e"),
   781 => (x"e3",x"c2",x"49",x"bf"),
   782 => (x"a1",x"c1",x"48",x"e8"),
   783 => (x"ff",x"e2",x"71",x"78"),
   784 => (x"c0",x"86",x"c4",x"87"),
   785 => (x"c2",x"48",x"cc",x"f7"),
   786 => (x"cc",x"78",x"f4",x"e3"),
   787 => (x"cc",x"f7",x"c0",x"87"),
   788 => (x"e0",x"c0",x"48",x"bf"),
   789 => (x"d0",x"f7",x"c0",x"80"),
   790 => (x"f0",x"e3",x"c2",x"58"),
   791 => (x"80",x"c1",x"48",x"bf"),
   792 => (x"58",x"f4",x"e3",x"c2"),
   793 => (x"00",x"0d",x"cc",x"27"),
   794 => (x"bf",x"97",x"bf",x"00"),
   795 => (x"c2",x"02",x"9d",x"4d"),
   796 => (x"e5",x"c3",x"87",x"e5"),
   797 => (x"de",x"c2",x"02",x"ad"),
   798 => (x"cc",x"f7",x"c0",x"87"),
   799 => (x"a3",x"cb",x"4b",x"bf"),
   800 => (x"cf",x"4c",x"11",x"49"),
   801 => (x"d2",x"c1",x"05",x"ac"),
   802 => (x"df",x"49",x"75",x"87"),
   803 => (x"cd",x"89",x"c1",x"99"),
   804 => (x"c4",x"ec",x"c2",x"91"),
   805 => (x"4a",x"a3",x"c1",x"81"),
   806 => (x"a3",x"c3",x"51",x"12"),
   807 => (x"c5",x"51",x"12",x"4a"),
   808 => (x"51",x"12",x"4a",x"a3"),
   809 => (x"12",x"4a",x"a3",x"c7"),
   810 => (x"4a",x"a3",x"c9",x"51"),
   811 => (x"a3",x"ce",x"51",x"12"),
   812 => (x"d0",x"51",x"12",x"4a"),
   813 => (x"51",x"12",x"4a",x"a3"),
   814 => (x"12",x"4a",x"a3",x"d2"),
   815 => (x"4a",x"a3",x"d4",x"51"),
   816 => (x"a3",x"d6",x"51",x"12"),
   817 => (x"d8",x"51",x"12",x"4a"),
   818 => (x"51",x"12",x"4a",x"a3"),
   819 => (x"12",x"4a",x"a3",x"dc"),
   820 => (x"4a",x"a3",x"de",x"51"),
   821 => (x"7e",x"c1",x"51",x"12"),
   822 => (x"74",x"87",x"fc",x"c0"),
   823 => (x"05",x"99",x"c8",x"49"),
   824 => (x"74",x"87",x"ed",x"c0"),
   825 => (x"05",x"99",x"d0",x"49"),
   826 => (x"e0",x"c0",x"87",x"d3"),
   827 => (x"cc",x"c0",x"02",x"66"),
   828 => (x"c0",x"49",x"73",x"87"),
   829 => (x"70",x"0f",x"66",x"e0"),
   830 => (x"d3",x"c0",x"02",x"98"),
   831 => (x"c0",x"05",x"6e",x"87"),
   832 => (x"ec",x"c2",x"87",x"c6"),
   833 => (x"50",x"c0",x"48",x"c4"),
   834 => (x"bf",x"cc",x"f7",x"c0"),
   835 => (x"87",x"e9",x"c2",x"48"),
   836 => (x"48",x"d1",x"ec",x"c2"),
   837 => (x"c2",x"7e",x"50",x"c0"),
   838 => (x"49",x"bf",x"c0",x"ec"),
   839 => (x"bf",x"f0",x"e3",x"c2"),
   840 => (x"04",x"aa",x"71",x"4a"),
   841 => (x"cf",x"87",x"f5",x"fb"),
   842 => (x"f8",x"ff",x"ff",x"ff"),
   843 => (x"e4",x"f0",x"c2",x"4c"),
   844 => (x"c8",x"c0",x"05",x"bf"),
   845 => (x"fc",x"eb",x"c2",x"87"),
   846 => (x"fa",x"c1",x"02",x"bf"),
   847 => (x"ec",x"e3",x"c2",x"87"),
   848 => (x"f9",x"ec",x"49",x"bf"),
   849 => (x"f0",x"e3",x"c2",x"87"),
   850 => (x"48",x"a6",x"c4",x"58"),
   851 => (x"bf",x"ec",x"e3",x"c2"),
   852 => (x"fc",x"eb",x"c2",x"78"),
   853 => (x"db",x"c0",x"02",x"bf"),
   854 => (x"49",x"66",x"c4",x"87"),
   855 => (x"a9",x"74",x"99",x"74"),
   856 => (x"87",x"c8",x"c0",x"02"),
   857 => (x"c0",x"48",x"a6",x"c8"),
   858 => (x"87",x"e7",x"c0",x"78"),
   859 => (x"c1",x"48",x"a6",x"c8"),
   860 => (x"87",x"df",x"c0",x"78"),
   861 => (x"cf",x"49",x"66",x"c4"),
   862 => (x"a9",x"99",x"f8",x"ff"),
   863 => (x"87",x"c8",x"c0",x"02"),
   864 => (x"c0",x"48",x"a6",x"cc"),
   865 => (x"87",x"c5",x"c0",x"78"),
   866 => (x"c1",x"48",x"a6",x"cc"),
   867 => (x"48",x"a6",x"c8",x"78"),
   868 => (x"c8",x"78",x"66",x"cc"),
   869 => (x"de",x"c0",x"05",x"66"),
   870 => (x"49",x"66",x"c4",x"87"),
   871 => (x"eb",x"c2",x"89",x"c2"),
   872 => (x"c2",x"91",x"bf",x"f4"),
   873 => (x"48",x"bf",x"d0",x"f0"),
   874 => (x"e3",x"c2",x"80",x"71"),
   875 => (x"e3",x"c2",x"58",x"ec"),
   876 => (x"78",x"c0",x"48",x"f0"),
   877 => (x"c0",x"87",x"d5",x"f9"),
   878 => (x"ff",x"ff",x"cf",x"48"),
   879 => (x"f0",x"4c",x"f8",x"ff"),
   880 => (x"26",x"4d",x"26",x"8e"),
   881 => (x"26",x"4b",x"26",x"4c"),
   882 => (x"00",x"00",x"00",x"4f"),
   883 => (x"00",x"00",x"00",x"00"),
   884 => (x"ff",x"ff",x"ff",x"ff"),
   885 => (x"00",x"00",x"0d",x"dc"),
   886 => (x"00",x"00",x"0d",x"e8"),
   887 => (x"33",x"54",x"41",x"46"),
   888 => (x"20",x"20",x"20",x"32"),
   889 => (x"00",x"00",x"00",x"00"),
   890 => (x"31",x"54",x"41",x"46"),
   891 => (x"20",x"20",x"20",x"36"),
   892 => (x"d4",x"ff",x"1e",x"00"),
   893 => (x"78",x"ff",x"c3",x"48"),
   894 => (x"4f",x"26",x"48",x"68"),
   895 => (x"48",x"d4",x"ff",x"1e"),
   896 => (x"ff",x"78",x"ff",x"c3"),
   897 => (x"e1",x"c0",x"48",x"d0"),
   898 => (x"48",x"d4",x"ff",x"78"),
   899 => (x"4f",x"26",x"78",x"d4"),
   900 => (x"48",x"d0",x"ff",x"1e"),
   901 => (x"26",x"78",x"e0",x"c0"),
   902 => (x"d4",x"ff",x"1e",x"4f"),
   903 => (x"99",x"49",x"70",x"87"),
   904 => (x"c0",x"87",x"c6",x"02"),
   905 => (x"f1",x"05",x"a9",x"fb"),
   906 => (x"26",x"48",x"71",x"87"),
   907 => (x"5b",x"5e",x"0e",x"4f"),
   908 => (x"4b",x"71",x"0e",x"5c"),
   909 => (x"f8",x"fe",x"4c",x"c0"),
   910 => (x"99",x"49",x"70",x"87"),
   911 => (x"87",x"f9",x"c0",x"02"),
   912 => (x"02",x"a9",x"ec",x"c0"),
   913 => (x"c0",x"87",x"f2",x"c0"),
   914 => (x"c0",x"02",x"a9",x"fb"),
   915 => (x"66",x"cc",x"87",x"eb"),
   916 => (x"c7",x"03",x"ac",x"b7"),
   917 => (x"02",x"66",x"d0",x"87"),
   918 => (x"53",x"71",x"87",x"c2"),
   919 => (x"c2",x"02",x"99",x"71"),
   920 => (x"fe",x"84",x"c1",x"87"),
   921 => (x"49",x"70",x"87",x"cb"),
   922 => (x"87",x"cd",x"02",x"99"),
   923 => (x"02",x"a9",x"ec",x"c0"),
   924 => (x"fb",x"c0",x"87",x"c7"),
   925 => (x"d5",x"ff",x"05",x"a9"),
   926 => (x"02",x"66",x"d0",x"87"),
   927 => (x"97",x"c0",x"87",x"c3"),
   928 => (x"a9",x"ec",x"c0",x"7b"),
   929 => (x"74",x"87",x"c4",x"05"),
   930 => (x"74",x"87",x"c5",x"4a"),
   931 => (x"8a",x"0a",x"c0",x"4a"),
   932 => (x"4c",x"26",x"48",x"72"),
   933 => (x"4f",x"26",x"4b",x"26"),
   934 => (x"87",x"d5",x"fd",x"1e"),
   935 => (x"c0",x"4a",x"49",x"70"),
   936 => (x"c9",x"04",x"aa",x"f0"),
   937 => (x"aa",x"f9",x"c0",x"87"),
   938 => (x"c0",x"87",x"c3",x"01"),
   939 => (x"c1",x"c1",x"8a",x"f0"),
   940 => (x"87",x"c9",x"04",x"aa"),
   941 => (x"01",x"aa",x"da",x"c1"),
   942 => (x"f7",x"c0",x"87",x"c3"),
   943 => (x"26",x"48",x"72",x"8a"),
   944 => (x"5b",x"5e",x"0e",x"4f"),
   945 => (x"f8",x"0e",x"5d",x"5c"),
   946 => (x"c0",x"4c",x"71",x"86"),
   947 => (x"87",x"ec",x"fc",x"7e"),
   948 => (x"fd",x"c0",x"4b",x"c0"),
   949 => (x"49",x"bf",x"97",x"e0"),
   950 => (x"cf",x"04",x"a9",x"c0"),
   951 => (x"87",x"f9",x"fc",x"87"),
   952 => (x"fd",x"c0",x"83",x"c1"),
   953 => (x"49",x"bf",x"97",x"e0"),
   954 => (x"87",x"f1",x"06",x"ab"),
   955 => (x"97",x"e0",x"fd",x"c0"),
   956 => (x"87",x"cf",x"02",x"bf"),
   957 => (x"70",x"87",x"fa",x"fb"),
   958 => (x"c6",x"02",x"99",x"49"),
   959 => (x"a9",x"ec",x"c0",x"87"),
   960 => (x"c0",x"87",x"f1",x"05"),
   961 => (x"87",x"e9",x"fb",x"4b"),
   962 => (x"e4",x"fb",x"4d",x"70"),
   963 => (x"58",x"a6",x"c8",x"87"),
   964 => (x"70",x"87",x"de",x"fb"),
   965 => (x"c8",x"83",x"c1",x"4a"),
   966 => (x"69",x"97",x"49",x"a4"),
   967 => (x"da",x"05",x"ad",x"49"),
   968 => (x"49",x"a4",x"c9",x"87"),
   969 => (x"c4",x"49",x"69",x"97"),
   970 => (x"ce",x"05",x"a9",x"66"),
   971 => (x"49",x"a4",x"ca",x"87"),
   972 => (x"aa",x"49",x"69",x"97"),
   973 => (x"c1",x"87",x"c4",x"05"),
   974 => (x"c0",x"87",x"d0",x"7e"),
   975 => (x"c6",x"02",x"ad",x"ec"),
   976 => (x"ad",x"fb",x"c0",x"87"),
   977 => (x"c0",x"87",x"c4",x"05"),
   978 => (x"6e",x"7e",x"c1",x"4b"),
   979 => (x"87",x"f5",x"fe",x"02"),
   980 => (x"73",x"87",x"fd",x"fa"),
   981 => (x"26",x"8e",x"f8",x"48"),
   982 => (x"26",x"4c",x"26",x"4d"),
   983 => (x"00",x"4f",x"26",x"4b"),
   984 => (x"1e",x"73",x"1e",x"00"),
   985 => (x"c8",x"4b",x"d4",x"ff"),
   986 => (x"d0",x"ff",x"4a",x"66"),
   987 => (x"78",x"c5",x"c8",x"48"),
   988 => (x"c1",x"48",x"d4",x"ff"),
   989 => (x"7b",x"11",x"78",x"d4"),
   990 => (x"f9",x"05",x"8a",x"c1"),
   991 => (x"48",x"d0",x"ff",x"87"),
   992 => (x"4b",x"26",x"78",x"c4"),
   993 => (x"5e",x"0e",x"4f",x"26"),
   994 => (x"0e",x"5d",x"5c",x"5b"),
   995 => (x"7e",x"71",x"86",x"f8"),
   996 => (x"f0",x"c2",x"1e",x"6e"),
   997 => (x"dc",x"e5",x"49",x"f4"),
   998 => (x"70",x"86",x"c4",x"87"),
   999 => (x"e4",x"c4",x"02",x"98"),
  1000 => (x"e4",x"ec",x"c1",x"87"),
  1001 => (x"49",x"6e",x"4c",x"bf"),
  1002 => (x"c8",x"87",x"d6",x"fc"),
  1003 => (x"98",x"70",x"58",x"a6"),
  1004 => (x"c4",x"87",x"c5",x"05"),
  1005 => (x"78",x"c1",x"48",x"a6"),
  1006 => (x"c5",x"48",x"d0",x"ff"),
  1007 => (x"48",x"d4",x"ff",x"78"),
  1008 => (x"c4",x"78",x"d5",x"c1"),
  1009 => (x"89",x"c1",x"49",x"66"),
  1010 => (x"ec",x"c1",x"31",x"c6"),
  1011 => (x"4a",x"bf",x"97",x"dc"),
  1012 => (x"ff",x"b0",x"71",x"48"),
  1013 => (x"ff",x"78",x"08",x"d4"),
  1014 => (x"78",x"c4",x"48",x"d0"),
  1015 => (x"97",x"f0",x"f0",x"c2"),
  1016 => (x"99",x"d0",x"49",x"bf"),
  1017 => (x"c5",x"87",x"dd",x"02"),
  1018 => (x"48",x"d4",x"ff",x"78"),
  1019 => (x"c0",x"78",x"d6",x"c1"),
  1020 => (x"48",x"d4",x"ff",x"4a"),
  1021 => (x"c1",x"78",x"ff",x"c3"),
  1022 => (x"aa",x"e0",x"c0",x"82"),
  1023 => (x"ff",x"87",x"f2",x"04"),
  1024 => (x"78",x"c4",x"48",x"d0"),
  1025 => (x"c3",x"48",x"d4",x"ff"),
  1026 => (x"d0",x"ff",x"78",x"ff"),
  1027 => (x"ff",x"78",x"c5",x"48"),
  1028 => (x"d3",x"c1",x"48",x"d4"),
  1029 => (x"ff",x"78",x"c1",x"78"),
  1030 => (x"78",x"c4",x"48",x"d0"),
  1031 => (x"06",x"ac",x"b7",x"c0"),
  1032 => (x"c2",x"87",x"cb",x"c2"),
  1033 => (x"4b",x"bf",x"fc",x"f0"),
  1034 => (x"73",x"7e",x"74",x"8c"),
  1035 => (x"dd",x"c1",x"02",x"9b"),
  1036 => (x"4d",x"c0",x"c8",x"87"),
  1037 => (x"ab",x"b7",x"c0",x"8b"),
  1038 => (x"c8",x"87",x"c6",x"03"),
  1039 => (x"c0",x"4d",x"a3",x"c0"),
  1040 => (x"f0",x"f0",x"c2",x"4b"),
  1041 => (x"d0",x"49",x"bf",x"97"),
  1042 => (x"87",x"cf",x"02",x"99"),
  1043 => (x"f0",x"c2",x"1e",x"c0"),
  1044 => (x"e1",x"e7",x"49",x"f4"),
  1045 => (x"70",x"86",x"c4",x"87"),
  1046 => (x"c2",x"87",x"d8",x"4c"),
  1047 => (x"c2",x"1e",x"f4",x"e3"),
  1048 => (x"e7",x"49",x"f4",x"f0"),
  1049 => (x"4c",x"70",x"87",x"d0"),
  1050 => (x"e3",x"c2",x"1e",x"75"),
  1051 => (x"f0",x"fb",x"49",x"f4"),
  1052 => (x"74",x"86",x"c8",x"87"),
  1053 => (x"87",x"c5",x"05",x"9c"),
  1054 => (x"ca",x"c1",x"48",x"c0"),
  1055 => (x"c2",x"1e",x"c1",x"87"),
  1056 => (x"e5",x"49",x"f4",x"f0"),
  1057 => (x"86",x"c4",x"87",x"d5"),
  1058 => (x"fe",x"05",x"9b",x"73"),
  1059 => (x"4c",x"6e",x"87",x"e3"),
  1060 => (x"06",x"ac",x"b7",x"c0"),
  1061 => (x"f0",x"c2",x"87",x"d1"),
  1062 => (x"78",x"c0",x"48",x"f4"),
  1063 => (x"78",x"c0",x"80",x"d0"),
  1064 => (x"f1",x"c2",x"80",x"f4"),
  1065 => (x"c0",x"78",x"bf",x"c0"),
  1066 => (x"fd",x"01",x"ac",x"b7"),
  1067 => (x"d0",x"ff",x"87",x"f5"),
  1068 => (x"ff",x"78",x"c5",x"48"),
  1069 => (x"d3",x"c1",x"48",x"d4"),
  1070 => (x"ff",x"78",x"c0",x"78"),
  1071 => (x"78",x"c4",x"48",x"d0"),
  1072 => (x"c2",x"c0",x"48",x"c1"),
  1073 => (x"f8",x"48",x"c0",x"87"),
  1074 => (x"26",x"4d",x"26",x"8e"),
  1075 => (x"26",x"4b",x"26",x"4c"),
  1076 => (x"5b",x"5e",x"0e",x"4f"),
  1077 => (x"fc",x"0e",x"5d",x"5c"),
  1078 => (x"c0",x"4d",x"71",x"86"),
  1079 => (x"04",x"ad",x"4c",x"4b"),
  1080 => (x"c0",x"87",x"e8",x"c0"),
  1081 => (x"74",x"1e",x"c1",x"fb"),
  1082 => (x"87",x"c4",x"02",x"9c"),
  1083 => (x"87",x"c2",x"4a",x"c0"),
  1084 => (x"49",x"72",x"4a",x"c1"),
  1085 => (x"c4",x"87",x"df",x"eb"),
  1086 => (x"c1",x"7e",x"70",x"86"),
  1087 => (x"c2",x"05",x"6e",x"83"),
  1088 => (x"c1",x"4b",x"75",x"87"),
  1089 => (x"06",x"ab",x"75",x"84"),
  1090 => (x"6e",x"87",x"d8",x"ff"),
  1091 => (x"26",x"8e",x"fc",x"48"),
  1092 => (x"26",x"4c",x"26",x"4d"),
  1093 => (x"0e",x"4f",x"26",x"4b"),
  1094 => (x"0e",x"5c",x"5b",x"5e"),
  1095 => (x"66",x"cc",x"4b",x"71"),
  1096 => (x"4c",x"87",x"d8",x"02"),
  1097 => (x"02",x"8c",x"f0",x"c0"),
  1098 => (x"4a",x"74",x"87",x"d8"),
  1099 => (x"d1",x"02",x"8a",x"c1"),
  1100 => (x"cd",x"02",x"8a",x"87"),
  1101 => (x"c9",x"02",x"8a",x"87"),
  1102 => (x"73",x"87",x"d9",x"87"),
  1103 => (x"87",x"c6",x"f9",x"49"),
  1104 => (x"1e",x"74",x"87",x"d2"),
  1105 => (x"da",x"c1",x"49",x"c0"),
  1106 => (x"1e",x"74",x"87",x"de"),
  1107 => (x"da",x"c1",x"49",x"73"),
  1108 => (x"86",x"c8",x"87",x"d6"),
  1109 => (x"4b",x"26",x"4c",x"26"),
  1110 => (x"5e",x"0e",x"4f",x"26"),
  1111 => (x"0e",x"5d",x"5c",x"5b"),
  1112 => (x"4c",x"71",x"86",x"fc"),
  1113 => (x"c2",x"91",x"de",x"49"),
  1114 => (x"71",x"4d",x"e0",x"f1"),
  1115 => (x"02",x"6d",x"97",x"85"),
  1116 => (x"c2",x"87",x"dc",x"c1"),
  1117 => (x"49",x"bf",x"d0",x"f1"),
  1118 => (x"fd",x"71",x"81",x"74"),
  1119 => (x"7e",x"70",x"87",x"d3"),
  1120 => (x"c0",x"02",x"98",x"48"),
  1121 => (x"f1",x"c2",x"87",x"f2"),
  1122 => (x"4a",x"70",x"4b",x"d4"),
  1123 => (x"fe",x"fe",x"49",x"cb"),
  1124 => (x"4b",x"74",x"87",x"d2"),
  1125 => (x"ec",x"c1",x"93",x"cc"),
  1126 => (x"83",x"c4",x"83",x"e8"),
  1127 => (x"7b",x"dc",x"c7",x"c1"),
  1128 => (x"c4",x"c1",x"49",x"74"),
  1129 => (x"7b",x"75",x"87",x"d6"),
  1130 => (x"97",x"e0",x"ec",x"c1"),
  1131 => (x"c2",x"1e",x"49",x"bf"),
  1132 => (x"fd",x"49",x"d4",x"f1"),
  1133 => (x"86",x"c4",x"87",x"e1"),
  1134 => (x"c3",x"c1",x"49",x"74"),
  1135 => (x"49",x"c0",x"87",x"fe"),
  1136 => (x"87",x"d9",x"c5",x"c1"),
  1137 => (x"48",x"ec",x"f0",x"c2"),
  1138 => (x"c0",x"49",x"50",x"c0"),
  1139 => (x"fc",x"87",x"c8",x"e2"),
  1140 => (x"26",x"4d",x"26",x"8e"),
  1141 => (x"26",x"4b",x"26",x"4c"),
  1142 => (x"00",x"00",x"00",x"4f"),
  1143 => (x"64",x"61",x"6f",x"4c"),
  1144 => (x"2e",x"67",x"6e",x"69"),
  1145 => (x"1e",x"00",x"2e",x"2e"),
  1146 => (x"4b",x"71",x"1e",x"73"),
  1147 => (x"d0",x"f1",x"c2",x"49"),
  1148 => (x"fb",x"71",x"81",x"bf"),
  1149 => (x"4a",x"70",x"87",x"db"),
  1150 => (x"87",x"c4",x"02",x"9a"),
  1151 => (x"87",x"dc",x"e6",x"49"),
  1152 => (x"48",x"d0",x"f1",x"c2"),
  1153 => (x"49",x"73",x"78",x"c0"),
  1154 => (x"26",x"87",x"fa",x"c1"),
  1155 => (x"1e",x"4f",x"26",x"4b"),
  1156 => (x"4b",x"71",x"1e",x"73"),
  1157 => (x"02",x"4a",x"a3",x"c4"),
  1158 => (x"c1",x"87",x"d0",x"c1"),
  1159 => (x"87",x"dc",x"02",x"8a"),
  1160 => (x"f2",x"c0",x"02",x"8a"),
  1161 => (x"c1",x"05",x"8a",x"87"),
  1162 => (x"f1",x"c2",x"87",x"d3"),
  1163 => (x"c1",x"02",x"bf",x"d0"),
  1164 => (x"c1",x"48",x"87",x"cb"),
  1165 => (x"d4",x"f1",x"c2",x"88"),
  1166 => (x"87",x"c1",x"c1",x"58"),
  1167 => (x"bf",x"d0",x"f1",x"c2"),
  1168 => (x"c2",x"89",x"c6",x"49"),
  1169 => (x"c0",x"59",x"d4",x"f1"),
  1170 => (x"c0",x"03",x"a9",x"b7"),
  1171 => (x"f1",x"c2",x"87",x"ef"),
  1172 => (x"78",x"c0",x"48",x"d0"),
  1173 => (x"c2",x"87",x"e6",x"c0"),
  1174 => (x"02",x"bf",x"cc",x"f1"),
  1175 => (x"f1",x"c2",x"87",x"df"),
  1176 => (x"c1",x"48",x"bf",x"d0"),
  1177 => (x"d4",x"f1",x"c2",x"80"),
  1178 => (x"c2",x"87",x"d2",x"58"),
  1179 => (x"02",x"bf",x"cc",x"f1"),
  1180 => (x"f1",x"c2",x"87",x"cb"),
  1181 => (x"c6",x"48",x"bf",x"d0"),
  1182 => (x"d4",x"f1",x"c2",x"80"),
  1183 => (x"c4",x"49",x"73",x"58"),
  1184 => (x"26",x"4b",x"26",x"87"),
  1185 => (x"5b",x"5e",x"0e",x"4f"),
  1186 => (x"f0",x"0e",x"5d",x"5c"),
  1187 => (x"59",x"a6",x"d0",x"86"),
  1188 => (x"4d",x"f4",x"e3",x"c2"),
  1189 => (x"f1",x"c2",x"4c",x"c0"),
  1190 => (x"78",x"c1",x"48",x"cc"),
  1191 => (x"c0",x"48",x"a6",x"c4"),
  1192 => (x"c2",x"7e",x"75",x"78"),
  1193 => (x"48",x"bf",x"d0",x"f1"),
  1194 => (x"c0",x"06",x"a8",x"c0"),
  1195 => (x"7e",x"75",x"87",x"fa"),
  1196 => (x"48",x"f4",x"e3",x"c2"),
  1197 => (x"ef",x"c0",x"02",x"98"),
  1198 => (x"c1",x"fb",x"c0",x"87"),
  1199 => (x"02",x"66",x"c8",x"1e"),
  1200 => (x"4d",x"c0",x"87",x"c4"),
  1201 => (x"4d",x"c1",x"87",x"c2"),
  1202 => (x"c9",x"e4",x"49",x"75"),
  1203 => (x"70",x"86",x"c4",x"87"),
  1204 => (x"c4",x"84",x"c1",x"7e"),
  1205 => (x"80",x"c1",x"48",x"66"),
  1206 => (x"c2",x"58",x"a6",x"c8"),
  1207 => (x"ac",x"bf",x"d0",x"f1"),
  1208 => (x"6e",x"87",x"c5",x"03"),
  1209 => (x"87",x"d1",x"ff",x"05"),
  1210 => (x"4c",x"c0",x"4d",x"6e"),
  1211 => (x"c3",x"02",x"9d",x"75"),
  1212 => (x"fb",x"c0",x"87",x"de"),
  1213 => (x"66",x"c8",x"1e",x"c1"),
  1214 => (x"cc",x"87",x"c7",x"02"),
  1215 => (x"78",x"c0",x"48",x"a6"),
  1216 => (x"a6",x"cc",x"87",x"c5"),
  1217 => (x"cc",x"78",x"c1",x"48"),
  1218 => (x"c9",x"e3",x"49",x"66"),
  1219 => (x"70",x"86",x"c4",x"87"),
  1220 => (x"02",x"98",x"48",x"7e"),
  1221 => (x"49",x"87",x"e6",x"c2"),
  1222 => (x"69",x"97",x"81",x"cb"),
  1223 => (x"02",x"99",x"d0",x"49"),
  1224 => (x"c1",x"87",x"d6",x"c1"),
  1225 => (x"74",x"4a",x"e7",x"c7"),
  1226 => (x"c1",x"91",x"cc",x"49"),
  1227 => (x"72",x"81",x"e8",x"ec"),
  1228 => (x"c3",x"81",x"c8",x"79"),
  1229 => (x"49",x"74",x"51",x"ff"),
  1230 => (x"f1",x"c2",x"91",x"de"),
  1231 => (x"85",x"71",x"4d",x"e0"),
  1232 => (x"7d",x"97",x"c1",x"c2"),
  1233 => (x"c0",x"49",x"a5",x"c1"),
  1234 => (x"ec",x"c2",x"51",x"e0"),
  1235 => (x"02",x"bf",x"97",x"c4"),
  1236 => (x"84",x"c1",x"87",x"d2"),
  1237 => (x"c2",x"4b",x"a5",x"c2"),
  1238 => (x"db",x"4a",x"c4",x"ec"),
  1239 => (x"c3",x"f7",x"fe",x"49"),
  1240 => (x"87",x"d9",x"c1",x"87"),
  1241 => (x"c0",x"49",x"a5",x"cd"),
  1242 => (x"c2",x"84",x"c1",x"51"),
  1243 => (x"4a",x"6e",x"4b",x"a5"),
  1244 => (x"f6",x"fe",x"49",x"cb"),
  1245 => (x"c4",x"c1",x"87",x"ee"),
  1246 => (x"cc",x"49",x"74",x"87"),
  1247 => (x"e8",x"ec",x"c1",x"91"),
  1248 => (x"da",x"c5",x"c1",x"81"),
  1249 => (x"c4",x"ec",x"c2",x"79"),
  1250 => (x"d8",x"02",x"bf",x"97"),
  1251 => (x"de",x"49",x"74",x"87"),
  1252 => (x"c2",x"84",x"c1",x"91"),
  1253 => (x"71",x"4b",x"e0",x"f1"),
  1254 => (x"c4",x"ec",x"c2",x"83"),
  1255 => (x"fe",x"49",x"dd",x"4a"),
  1256 => (x"d8",x"87",x"c1",x"f6"),
  1257 => (x"de",x"4b",x"74",x"87"),
  1258 => (x"e0",x"f1",x"c2",x"93"),
  1259 => (x"49",x"a3",x"cb",x"83"),
  1260 => (x"84",x"c1",x"51",x"c0"),
  1261 => (x"cb",x"4a",x"6e",x"73"),
  1262 => (x"e7",x"f5",x"fe",x"49"),
  1263 => (x"48",x"66",x"c4",x"87"),
  1264 => (x"a6",x"c8",x"80",x"c1"),
  1265 => (x"03",x"ac",x"c7",x"58"),
  1266 => (x"6e",x"87",x"c5",x"c0"),
  1267 => (x"87",x"e2",x"fc",x"05"),
  1268 => (x"c0",x"03",x"ac",x"c7"),
  1269 => (x"f1",x"c2",x"87",x"e6"),
  1270 => (x"78",x"c0",x"48",x"cc"),
  1271 => (x"4a",x"da",x"c5",x"c1"),
  1272 => (x"91",x"cc",x"49",x"74"),
  1273 => (x"81",x"e8",x"ec",x"c1"),
  1274 => (x"49",x"74",x"79",x"72"),
  1275 => (x"f1",x"c2",x"91",x"de"),
  1276 => (x"51",x"c0",x"81",x"e0"),
  1277 => (x"ac",x"c7",x"84",x"c1"),
  1278 => (x"87",x"da",x"ff",x"04"),
  1279 => (x"48",x"c4",x"ee",x"c1"),
  1280 => (x"80",x"f7",x"50",x"c0"),
  1281 => (x"40",x"f1",x"d1",x"c1"),
  1282 => (x"78",x"e4",x"d0",x"c1"),
  1283 => (x"c8",x"c1",x"80",x"c8"),
  1284 => (x"66",x"cc",x"78",x"cf"),
  1285 => (x"e3",x"fa",x"c0",x"49"),
  1286 => (x"26",x"8e",x"f0",x"87"),
  1287 => (x"26",x"4c",x"26",x"4d"),
  1288 => (x"00",x"4f",x"26",x"4b"),
  1289 => (x"61",x"42",x"20",x"80"),
  1290 => (x"1e",x"00",x"6b",x"63"),
  1291 => (x"4b",x"71",x"1e",x"73"),
  1292 => (x"c1",x"91",x"cc",x"49"),
  1293 => (x"c8",x"81",x"e8",x"ec"),
  1294 => (x"ec",x"c1",x"4a",x"a1"),
  1295 => (x"50",x"12",x"48",x"dc"),
  1296 => (x"c0",x"4a",x"a1",x"c9"),
  1297 => (x"12",x"48",x"e0",x"fd"),
  1298 => (x"c1",x"81",x"ca",x"50"),
  1299 => (x"11",x"48",x"e0",x"ec"),
  1300 => (x"e0",x"ec",x"c1",x"50"),
  1301 => (x"1e",x"49",x"bf",x"97"),
  1302 => (x"fa",x"f2",x"49",x"c0"),
  1303 => (x"f8",x"49",x"73",x"87"),
  1304 => (x"8e",x"fc",x"87",x"e3"),
  1305 => (x"4f",x"26",x"4b",x"26"),
  1306 => (x"c0",x"49",x"c0",x"1e"),
  1307 => (x"26",x"87",x"ee",x"fa"),
  1308 => (x"4a",x"71",x"1e",x"4f"),
  1309 => (x"c1",x"91",x"cc",x"49"),
  1310 => (x"c8",x"81",x"e8",x"ec"),
  1311 => (x"ec",x"f0",x"c2",x"81"),
  1312 => (x"c0",x"50",x"11",x"48"),
  1313 => (x"fe",x"49",x"a2",x"f0"),
  1314 => (x"c0",x"87",x"c1",x"f0"),
  1315 => (x"87",x"c7",x"d7",x"49"),
  1316 => (x"ff",x"1e",x"4f",x"26"),
  1317 => (x"ff",x"c3",x"4a",x"d4"),
  1318 => (x"48",x"d0",x"ff",x"7a"),
  1319 => (x"de",x"78",x"e1",x"c0"),
  1320 => (x"48",x"7a",x"71",x"7a"),
  1321 => (x"70",x"28",x"b7",x"c8"),
  1322 => (x"d0",x"48",x"71",x"7a"),
  1323 => (x"7a",x"70",x"28",x"b7"),
  1324 => (x"b7",x"d8",x"48",x"71"),
  1325 => (x"ff",x"7a",x"70",x"28"),
  1326 => (x"e0",x"c0",x"48",x"d0"),
  1327 => (x"0e",x"4f",x"26",x"78"),
  1328 => (x"5d",x"5c",x"5b",x"5e"),
  1329 => (x"71",x"86",x"f4",x"0e"),
  1330 => (x"91",x"cc",x"49",x"4d"),
  1331 => (x"81",x"e8",x"ec",x"c1"),
  1332 => (x"ca",x"4a",x"a1",x"c8"),
  1333 => (x"a6",x"c4",x"7e",x"a1"),
  1334 => (x"e8",x"f0",x"c2",x"48"),
  1335 => (x"97",x"6e",x"78",x"bf"),
  1336 => (x"66",x"c4",x"4b",x"bf"),
  1337 => (x"12",x"2c",x"73",x"4c"),
  1338 => (x"58",x"a6",x"cc",x"48"),
  1339 => (x"84",x"c1",x"9c",x"70"),
  1340 => (x"69",x"97",x"81",x"c9"),
  1341 => (x"04",x"ac",x"b7",x"49"),
  1342 => (x"4c",x"c0",x"87",x"c2"),
  1343 => (x"4a",x"bf",x"97",x"6e"),
  1344 => (x"72",x"49",x"66",x"c8"),
  1345 => (x"c4",x"b9",x"ff",x"31"),
  1346 => (x"48",x"74",x"99",x"66"),
  1347 => (x"4a",x"70",x"30",x"72"),
  1348 => (x"ec",x"f0",x"c2",x"b1"),
  1349 => (x"f9",x"fd",x"71",x"59"),
  1350 => (x"c2",x"1e",x"c7",x"87"),
  1351 => (x"1e",x"bf",x"c8",x"f1"),
  1352 => (x"1e",x"e8",x"ec",x"c1"),
  1353 => (x"97",x"ec",x"f0",x"c2"),
  1354 => (x"f4",x"c1",x"49",x"bf"),
  1355 => (x"c0",x"49",x"75",x"87"),
  1356 => (x"e8",x"87",x"c9",x"f6"),
  1357 => (x"26",x"4d",x"26",x"8e"),
  1358 => (x"26",x"4b",x"26",x"4c"),
  1359 => (x"1e",x"73",x"1e",x"4f"),
  1360 => (x"fd",x"49",x"4b",x"71"),
  1361 => (x"49",x"73",x"87",x"f9"),
  1362 => (x"26",x"87",x"f4",x"fd"),
  1363 => (x"1e",x"4f",x"26",x"4b"),
  1364 => (x"4b",x"71",x"1e",x"73"),
  1365 => (x"02",x"4a",x"a3",x"c2"),
  1366 => (x"8a",x"c1",x"87",x"d6"),
  1367 => (x"87",x"e2",x"c0",x"05"),
  1368 => (x"bf",x"c8",x"f1",x"c2"),
  1369 => (x"48",x"87",x"db",x"02"),
  1370 => (x"f1",x"c2",x"88",x"c1"),
  1371 => (x"87",x"d2",x"58",x"cc"),
  1372 => (x"bf",x"cc",x"f1",x"c2"),
  1373 => (x"c2",x"87",x"cb",x"02"),
  1374 => (x"48",x"bf",x"c8",x"f1"),
  1375 => (x"f1",x"c2",x"80",x"c1"),
  1376 => (x"1e",x"c7",x"58",x"cc"),
  1377 => (x"bf",x"c8",x"f1",x"c2"),
  1378 => (x"e8",x"ec",x"c1",x"1e"),
  1379 => (x"ec",x"f0",x"c2",x"1e"),
  1380 => (x"cc",x"49",x"bf",x"97"),
  1381 => (x"c0",x"49",x"73",x"87"),
  1382 => (x"f4",x"87",x"e1",x"f4"),
  1383 => (x"26",x"4b",x"26",x"8e"),
  1384 => (x"5b",x"5e",x"0e",x"4f"),
  1385 => (x"ff",x"0e",x"5d",x"5c"),
  1386 => (x"e4",x"c0",x"86",x"cc"),
  1387 => (x"a6",x"cc",x"59",x"a6"),
  1388 => (x"c4",x"78",x"c0",x"48"),
  1389 => (x"c4",x"78",x"c0",x"80"),
  1390 => (x"66",x"c8",x"c1",x"80"),
  1391 => (x"c1",x"80",x"c4",x"78"),
  1392 => (x"c1",x"80",x"c4",x"78"),
  1393 => (x"cc",x"f1",x"c2",x"78"),
  1394 => (x"e0",x"78",x"c1",x"48"),
  1395 => (x"c8",x"e1",x"87",x"ee"),
  1396 => (x"87",x"dd",x"e0",x"87"),
  1397 => (x"fb",x"c0",x"4c",x"70"),
  1398 => (x"f3",x"c1",x"02",x"ac"),
  1399 => (x"66",x"e0",x"c0",x"87"),
  1400 => (x"87",x"e8",x"c1",x"05"),
  1401 => (x"4a",x"66",x"c4",x"c1"),
  1402 => (x"7e",x"6a",x"82",x"c4"),
  1403 => (x"48",x"f8",x"e8",x"c1"),
  1404 => (x"41",x"20",x"49",x"6e"),
  1405 => (x"51",x"10",x"41",x"20"),
  1406 => (x"48",x"66",x"c4",x"c1"),
  1407 => (x"78",x"eb",x"d0",x"c1"),
  1408 => (x"81",x"c7",x"49",x"6a"),
  1409 => (x"c4",x"c1",x"51",x"74"),
  1410 => (x"81",x"c8",x"49",x"66"),
  1411 => (x"a6",x"d8",x"51",x"c1"),
  1412 => (x"c1",x"78",x"c2",x"48"),
  1413 => (x"c9",x"49",x"66",x"c4"),
  1414 => (x"c1",x"51",x"c0",x"81"),
  1415 => (x"ca",x"49",x"66",x"c4"),
  1416 => (x"c1",x"51",x"c0",x"81"),
  1417 => (x"6a",x"1e",x"d8",x"1e"),
  1418 => (x"ff",x"81",x"c8",x"49"),
  1419 => (x"c8",x"87",x"fe",x"df"),
  1420 => (x"66",x"c8",x"c1",x"86"),
  1421 => (x"01",x"a8",x"c0",x"48"),
  1422 => (x"a6",x"d0",x"87",x"c7"),
  1423 => (x"cf",x"78",x"c1",x"48"),
  1424 => (x"66",x"c8",x"c1",x"87"),
  1425 => (x"d8",x"88",x"c1",x"48"),
  1426 => (x"87",x"c4",x"58",x"a6"),
  1427 => (x"87",x"c9",x"df",x"ff"),
  1428 => (x"cd",x"02",x"9c",x"74"),
  1429 => (x"66",x"d0",x"87",x"d9"),
  1430 => (x"66",x"cc",x"c1",x"48"),
  1431 => (x"ce",x"cd",x"03",x"a8"),
  1432 => (x"48",x"a6",x"c8",x"87"),
  1433 => (x"ff",x"7e",x"78",x"c0"),
  1434 => (x"70",x"87",x"c6",x"de"),
  1435 => (x"ac",x"d0",x"c1",x"4c"),
  1436 => (x"87",x"e7",x"c2",x"05"),
  1437 => (x"6e",x"48",x"a6",x"c4"),
  1438 => (x"87",x"dc",x"e0",x"78"),
  1439 => (x"cc",x"48",x"7e",x"70"),
  1440 => (x"c5",x"06",x"a8",x"66"),
  1441 => (x"48",x"a6",x"cc",x"87"),
  1442 => (x"dd",x"ff",x"78",x"6e"),
  1443 => (x"4c",x"70",x"87",x"e3"),
  1444 => (x"05",x"ac",x"ec",x"c0"),
  1445 => (x"d0",x"87",x"ee",x"c1"),
  1446 => (x"91",x"cc",x"49",x"66"),
  1447 => (x"81",x"66",x"c4",x"c1"),
  1448 => (x"6a",x"4a",x"a1",x"c4"),
  1449 => (x"4a",x"a1",x"c8",x"4d"),
  1450 => (x"d1",x"c1",x"52",x"6e"),
  1451 => (x"dc",x"ff",x"79",x"f1"),
  1452 => (x"4c",x"70",x"87",x"ff"),
  1453 => (x"87",x"d9",x"02",x"9c"),
  1454 => (x"02",x"ac",x"fb",x"c0"),
  1455 => (x"55",x"74",x"87",x"d3"),
  1456 => (x"87",x"ed",x"dc",x"ff"),
  1457 => (x"02",x"9c",x"4c",x"70"),
  1458 => (x"fb",x"c0",x"87",x"c7"),
  1459 => (x"ed",x"ff",x"05",x"ac"),
  1460 => (x"55",x"e0",x"c0",x"87"),
  1461 => (x"c0",x"55",x"c1",x"c2"),
  1462 => (x"e0",x"c0",x"7d",x"97"),
  1463 => (x"66",x"c4",x"48",x"66"),
  1464 => (x"87",x"db",x"05",x"a8"),
  1465 => (x"d4",x"48",x"66",x"d0"),
  1466 => (x"ca",x"04",x"a8",x"66"),
  1467 => (x"48",x"66",x"d0",x"87"),
  1468 => (x"a6",x"d4",x"80",x"c1"),
  1469 => (x"d4",x"87",x"c8",x"58"),
  1470 => (x"88",x"c1",x"48",x"66"),
  1471 => (x"ff",x"58",x"a6",x"d8"),
  1472 => (x"70",x"87",x"ee",x"db"),
  1473 => (x"ac",x"d0",x"c1",x"4c"),
  1474 => (x"dc",x"87",x"c9",x"05"),
  1475 => (x"80",x"c1",x"48",x"66"),
  1476 => (x"58",x"a6",x"e0",x"c0"),
  1477 => (x"02",x"ac",x"d0",x"c1"),
  1478 => (x"6e",x"87",x"d9",x"fd"),
  1479 => (x"66",x"e0",x"c0",x"48"),
  1480 => (x"ea",x"c9",x"05",x"a8"),
  1481 => (x"a6",x"e4",x"c0",x"87"),
  1482 => (x"74",x"78",x"c0",x"48"),
  1483 => (x"88",x"fb",x"c0",x"48"),
  1484 => (x"70",x"58",x"a6",x"c8"),
  1485 => (x"dc",x"c9",x"02",x"98"),
  1486 => (x"88",x"cb",x"48",x"87"),
  1487 => (x"70",x"58",x"a6",x"c8"),
  1488 => (x"ce",x"c1",x"02",x"98"),
  1489 => (x"88",x"c9",x"48",x"87"),
  1490 => (x"70",x"58",x"a6",x"c8"),
  1491 => (x"fe",x"c3",x"02",x"98"),
  1492 => (x"88",x"c4",x"48",x"87"),
  1493 => (x"70",x"58",x"a6",x"c8"),
  1494 => (x"87",x"cf",x"02",x"98"),
  1495 => (x"c8",x"88",x"c1",x"48"),
  1496 => (x"98",x"70",x"58",x"a6"),
  1497 => (x"87",x"e7",x"c3",x"02"),
  1498 => (x"c8",x"87",x"db",x"c8"),
  1499 => (x"f0",x"c0",x"48",x"a6"),
  1500 => (x"fc",x"d9",x"ff",x"78"),
  1501 => (x"c0",x"4c",x"70",x"87"),
  1502 => (x"c3",x"02",x"ac",x"ec"),
  1503 => (x"5c",x"a6",x"cc",x"87"),
  1504 => (x"02",x"ac",x"ec",x"c0"),
  1505 => (x"d9",x"ff",x"87",x"cd"),
  1506 => (x"4c",x"70",x"87",x"e7"),
  1507 => (x"05",x"ac",x"ec",x"c0"),
  1508 => (x"c0",x"87",x"f3",x"ff"),
  1509 => (x"c0",x"02",x"ac",x"ec"),
  1510 => (x"d9",x"ff",x"87",x"c4"),
  1511 => (x"1e",x"c0",x"87",x"d3"),
  1512 => (x"66",x"d8",x"1e",x"ca"),
  1513 => (x"c1",x"91",x"cc",x"49"),
  1514 => (x"71",x"48",x"66",x"cc"),
  1515 => (x"58",x"a6",x"cc",x"80"),
  1516 => (x"c4",x"48",x"66",x"c8"),
  1517 => (x"58",x"a6",x"d0",x"80"),
  1518 => (x"49",x"bf",x"66",x"cc"),
  1519 => (x"87",x"ed",x"d9",x"ff"),
  1520 => (x"1e",x"de",x"1e",x"c1"),
  1521 => (x"49",x"bf",x"66",x"d4"),
  1522 => (x"87",x"e1",x"d9",x"ff"),
  1523 => (x"49",x"70",x"86",x"d0"),
  1524 => (x"88",x"08",x"c0",x"48"),
  1525 => (x"58",x"a6",x"ec",x"c0"),
  1526 => (x"c0",x"06",x"a8",x"c0"),
  1527 => (x"e8",x"c0",x"87",x"ee"),
  1528 => (x"a8",x"dd",x"48",x"66"),
  1529 => (x"87",x"e4",x"c0",x"03"),
  1530 => (x"49",x"bf",x"66",x"c4"),
  1531 => (x"81",x"66",x"e8",x"c0"),
  1532 => (x"c0",x"51",x"e0",x"c0"),
  1533 => (x"c1",x"49",x"66",x"e8"),
  1534 => (x"bf",x"66",x"c4",x"81"),
  1535 => (x"51",x"c1",x"c2",x"81"),
  1536 => (x"49",x"66",x"e8",x"c0"),
  1537 => (x"66",x"c4",x"81",x"c2"),
  1538 => (x"51",x"c0",x"81",x"bf"),
  1539 => (x"d0",x"c1",x"48",x"6e"),
  1540 => (x"49",x"6e",x"78",x"eb"),
  1541 => (x"66",x"d8",x"81",x"c8"),
  1542 => (x"c9",x"49",x"6e",x"51"),
  1543 => (x"51",x"66",x"dc",x"81"),
  1544 => (x"81",x"ca",x"49",x"6e"),
  1545 => (x"d8",x"51",x"66",x"c8"),
  1546 => (x"80",x"c1",x"48",x"66"),
  1547 => (x"d0",x"58",x"a6",x"dc"),
  1548 => (x"66",x"d4",x"48",x"66"),
  1549 => (x"cb",x"c0",x"04",x"a8"),
  1550 => (x"48",x"66",x"d0",x"87"),
  1551 => (x"a6",x"d4",x"80",x"c1"),
  1552 => (x"87",x"d1",x"c5",x"58"),
  1553 => (x"c1",x"48",x"66",x"d4"),
  1554 => (x"58",x"a6",x"d8",x"88"),
  1555 => (x"ff",x"87",x"c6",x"c5"),
  1556 => (x"c0",x"87",x"c5",x"d9"),
  1557 => (x"ff",x"58",x"a6",x"ec"),
  1558 => (x"c0",x"87",x"fd",x"d8"),
  1559 => (x"c0",x"58",x"a6",x"f0"),
  1560 => (x"c0",x"05",x"a8",x"ec"),
  1561 => (x"48",x"a6",x"87",x"c9"),
  1562 => (x"78",x"66",x"e8",x"c0"),
  1563 => (x"ff",x"87",x"c4",x"c0"),
  1564 => (x"d0",x"87",x"fe",x"d5"),
  1565 => (x"91",x"cc",x"49",x"66"),
  1566 => (x"48",x"66",x"c4",x"c1"),
  1567 => (x"a6",x"c8",x"80",x"71"),
  1568 => (x"4a",x"66",x"c4",x"58"),
  1569 => (x"66",x"c4",x"82",x"c8"),
  1570 => (x"c0",x"81",x"ca",x"49"),
  1571 => (x"c0",x"51",x"66",x"e8"),
  1572 => (x"c1",x"49",x"66",x"ec"),
  1573 => (x"66",x"e8",x"c0",x"81"),
  1574 => (x"71",x"48",x"c1",x"89"),
  1575 => (x"c1",x"49",x"70",x"30"),
  1576 => (x"7a",x"97",x"71",x"89"),
  1577 => (x"bf",x"e8",x"f0",x"c2"),
  1578 => (x"66",x"e8",x"c0",x"49"),
  1579 => (x"4a",x"6a",x"97",x"29"),
  1580 => (x"c0",x"98",x"71",x"48"),
  1581 => (x"c4",x"58",x"a6",x"f4"),
  1582 => (x"80",x"c4",x"48",x"66"),
  1583 => (x"c8",x"58",x"a6",x"cc"),
  1584 => (x"c0",x"4d",x"bf",x"66"),
  1585 => (x"6e",x"48",x"66",x"e0"),
  1586 => (x"c5",x"c0",x"02",x"a8"),
  1587 => (x"c0",x"7e",x"c0",x"87"),
  1588 => (x"7e",x"c1",x"87",x"c2"),
  1589 => (x"e0",x"c0",x"1e",x"6e"),
  1590 => (x"ff",x"49",x"75",x"1e"),
  1591 => (x"c8",x"87",x"ce",x"d5"),
  1592 => (x"c0",x"4c",x"70",x"86"),
  1593 => (x"c1",x"06",x"ac",x"b7"),
  1594 => (x"85",x"74",x"87",x"d4"),
  1595 => (x"49",x"bf",x"66",x"c8"),
  1596 => (x"75",x"81",x"e0",x"c0"),
  1597 => (x"e9",x"c1",x"4b",x"89"),
  1598 => (x"fe",x"71",x"4a",x"c4"),
  1599 => (x"c2",x"87",x"e5",x"e0"),
  1600 => (x"c0",x"7e",x"75",x"85"),
  1601 => (x"c1",x"48",x"66",x"e4"),
  1602 => (x"a6",x"e8",x"c0",x"80"),
  1603 => (x"66",x"f0",x"c0",x"58"),
  1604 => (x"70",x"81",x"c1",x"49"),
  1605 => (x"c5",x"c0",x"02",x"a9"),
  1606 => (x"c0",x"4d",x"c0",x"87"),
  1607 => (x"4d",x"c1",x"87",x"c2"),
  1608 => (x"66",x"cc",x"1e",x"75"),
  1609 => (x"e0",x"c0",x"49",x"bf"),
  1610 => (x"89",x"66",x"c4",x"81"),
  1611 => (x"66",x"c8",x"1e",x"71"),
  1612 => (x"f8",x"d3",x"ff",x"49"),
  1613 => (x"c0",x"86",x"c8",x"87"),
  1614 => (x"ff",x"01",x"a8",x"b7"),
  1615 => (x"e4",x"c0",x"87",x"c5"),
  1616 => (x"d3",x"c0",x"02",x"66"),
  1617 => (x"49",x"66",x"c4",x"87"),
  1618 => (x"e4",x"c0",x"81",x"c9"),
  1619 => (x"66",x"c4",x"51",x"66"),
  1620 => (x"ff",x"d2",x"c1",x"48"),
  1621 => (x"87",x"ce",x"c0",x"78"),
  1622 => (x"c9",x"49",x"66",x"c4"),
  1623 => (x"c4",x"51",x"c2",x"81"),
  1624 => (x"d4",x"c1",x"48",x"66"),
  1625 => (x"66",x"d0",x"78",x"fd"),
  1626 => (x"a8",x"66",x"d4",x"48"),
  1627 => (x"87",x"cb",x"c0",x"04"),
  1628 => (x"c1",x"48",x"66",x"d0"),
  1629 => (x"58",x"a6",x"d4",x"80"),
  1630 => (x"d4",x"87",x"da",x"c0"),
  1631 => (x"88",x"c1",x"48",x"66"),
  1632 => (x"c0",x"58",x"a6",x"d8"),
  1633 => (x"d2",x"ff",x"87",x"cf"),
  1634 => (x"4c",x"70",x"87",x"cf"),
  1635 => (x"ff",x"87",x"c6",x"c0"),
  1636 => (x"70",x"87",x"c6",x"d2"),
  1637 => (x"48",x"66",x"dc",x"4c"),
  1638 => (x"e0",x"c0",x"80",x"c1"),
  1639 => (x"9c",x"74",x"58",x"a6"),
  1640 => (x"87",x"cb",x"c0",x"02"),
  1641 => (x"c1",x"48",x"66",x"d0"),
  1642 => (x"04",x"a8",x"66",x"cc"),
  1643 => (x"d0",x"87",x"f2",x"f2"),
  1644 => (x"a8",x"c7",x"48",x"66"),
  1645 => (x"87",x"e1",x"c0",x"03"),
  1646 => (x"c2",x"4c",x"66",x"d0"),
  1647 => (x"c0",x"48",x"cc",x"f1"),
  1648 => (x"cc",x"49",x"74",x"78"),
  1649 => (x"66",x"c4",x"c1",x"91"),
  1650 => (x"4a",x"a1",x"c4",x"81"),
  1651 => (x"52",x"c0",x"4a",x"6a"),
  1652 => (x"c7",x"84",x"c1",x"79"),
  1653 => (x"e2",x"ff",x"04",x"ac"),
  1654 => (x"66",x"e0",x"c0",x"87"),
  1655 => (x"87",x"e2",x"c0",x"02"),
  1656 => (x"49",x"66",x"c4",x"c1"),
  1657 => (x"c1",x"81",x"d4",x"c1"),
  1658 => (x"c1",x"4a",x"66",x"c4"),
  1659 => (x"52",x"c0",x"82",x"dc"),
  1660 => (x"79",x"f1",x"d1",x"c1"),
  1661 => (x"49",x"66",x"c4",x"c1"),
  1662 => (x"c1",x"81",x"d8",x"c1"),
  1663 => (x"c0",x"79",x"c8",x"e9"),
  1664 => (x"c4",x"c1",x"87",x"d6"),
  1665 => (x"d4",x"c1",x"49",x"66"),
  1666 => (x"66",x"c4",x"c1",x"81"),
  1667 => (x"82",x"d8",x"c1",x"4a"),
  1668 => (x"7a",x"d0",x"e9",x"c1"),
  1669 => (x"79",x"e8",x"d1",x"c1"),
  1670 => (x"49",x"66",x"c4",x"c1"),
  1671 => (x"c1",x"81",x"e0",x"c1"),
  1672 => (x"ff",x"79",x"cf",x"d5"),
  1673 => (x"cc",x"87",x"e9",x"cf"),
  1674 => (x"cc",x"ff",x"48",x"66"),
  1675 => (x"26",x"4d",x"26",x"8e"),
  1676 => (x"26",x"4b",x"26",x"4c"),
  1677 => (x"00",x"00",x"00",x"4f"),
  1678 => (x"64",x"61",x"6f",x"4c"),
  1679 => (x"20",x"2e",x"2a",x"20"),
  1680 => (x"00",x"00",x"00",x"00"),
  1681 => (x"00",x"00",x"20",x"3a"),
  1682 => (x"61",x"42",x"20",x"80"),
  1683 => (x"00",x"00",x"6b",x"63"),
  1684 => (x"78",x"45",x"20",x"80"),
  1685 => (x"1e",x"00",x"74",x"69"),
  1686 => (x"f1",x"c2",x"1e",x"c7"),
  1687 => (x"c1",x"1e",x"bf",x"c8"),
  1688 => (x"c2",x"1e",x"e8",x"ec"),
  1689 => (x"bf",x"97",x"ec",x"f0"),
  1690 => (x"87",x"f5",x"ec",x"49"),
  1691 => (x"49",x"e8",x"ec",x"c1"),
  1692 => (x"87",x"d6",x"e2",x"c0"),
  1693 => (x"4f",x"26",x"8e",x"f4"),
  1694 => (x"c8",x"1e",x"73",x"1e"),
  1695 => (x"ee",x"c1",x"87",x"c3"),
  1696 => (x"ec",x"c1",x"48",x"c0"),
  1697 => (x"e8",x"fe",x"78",x"c8"),
  1698 => (x"e1",x"c0",x"49",x"a0"),
  1699 => (x"49",x"c7",x"87",x"fc"),
  1700 => (x"87",x"e8",x"e0",x"c0"),
  1701 => (x"e2",x"c0",x"49",x"c1"),
  1702 => (x"d4",x"ff",x"87",x"c3"),
  1703 => (x"78",x"ff",x"c3",x"48"),
  1704 => (x"48",x"d4",x"f1",x"c2"),
  1705 => (x"e3",x"fe",x"50",x"c0"),
  1706 => (x"98",x"70",x"87",x"e2"),
  1707 => (x"fe",x"87",x"cd",x"02"),
  1708 => (x"70",x"87",x"de",x"ed"),
  1709 => (x"87",x"c4",x"02",x"98"),
  1710 => (x"87",x"c2",x"4a",x"c1"),
  1711 => (x"9a",x"72",x"4a",x"c0"),
  1712 => (x"c1",x"87",x"c8",x"02"),
  1713 => (x"fe",x"49",x"d4",x"ec"),
  1714 => (x"c2",x"87",x"dc",x"d7"),
  1715 => (x"c0",x"48",x"c8",x"f1"),
  1716 => (x"ec",x"f0",x"c2",x"78"),
  1717 => (x"49",x"50",x"c0",x"48"),
  1718 => (x"c0",x"87",x"fc",x"fd"),
  1719 => (x"70",x"87",x"cd",x"f6"),
  1720 => (x"cb",x"02",x"9b",x"4b"),
  1721 => (x"c4",x"ee",x"c1",x"87"),
  1722 => (x"df",x"49",x"c7",x"5b"),
  1723 => (x"87",x"c6",x"87",x"ce"),
  1724 => (x"e0",x"c0",x"49",x"c0"),
  1725 => (x"c2",x"c3",x"87",x"e7"),
  1726 => (x"c8",x"e2",x"c0",x"87"),
  1727 => (x"d4",x"f0",x"c0",x"87"),
  1728 => (x"87",x"f5",x"ff",x"87"),
  1729 => (x"4f",x"26",x"4b",x"26"),
  1730 => (x"74",x"6f",x"6f",x"42"),
  1731 => (x"2e",x"67",x"6e",x"69"),
  1732 => (x"00",x"00",x"2e",x"2e"),
  1733 => (x"4f",x"20",x"44",x"53"),
  1734 => (x"00",x"00",x"00",x"4b"),
  1735 => (x"00",x"00",x"00",x"00"),
  1736 => (x"00",x"00",x"00",x"00"),
  1737 => (x"00",x"00",x"00",x"01"),
  1738 => (x"00",x"00",x"11",x"5a"),
  1739 => (x"00",x"00",x"2c",x"60"),
  1740 => (x"00",x"00",x"00",x"00"),
  1741 => (x"00",x"00",x"11",x"5a"),
  1742 => (x"00",x"00",x"2c",x"7e"),
  1743 => (x"00",x"00",x"00",x"00"),
  1744 => (x"00",x"00",x"11",x"5a"),
  1745 => (x"00",x"00",x"2c",x"9c"),
  1746 => (x"00",x"00",x"00",x"00"),
  1747 => (x"00",x"00",x"11",x"5a"),
  1748 => (x"00",x"00",x"2c",x"ba"),
  1749 => (x"00",x"00",x"00",x"00"),
  1750 => (x"00",x"00",x"11",x"5a"),
  1751 => (x"00",x"00",x"2c",x"d8"),
  1752 => (x"00",x"00",x"00",x"00"),
  1753 => (x"00",x"00",x"11",x"5a"),
  1754 => (x"00",x"00",x"2c",x"f6"),
  1755 => (x"00",x"00",x"00",x"00"),
  1756 => (x"00",x"00",x"11",x"5a"),
  1757 => (x"00",x"00",x"2d",x"14"),
  1758 => (x"00",x"00",x"00",x"00"),
  1759 => (x"00",x"00",x"14",x"71"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"12",x"0f"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"db",x"86",x"fc",x"1e"),
  1766 => (x"fc",x"7e",x"70",x"87"),
  1767 => (x"1e",x"4f",x"26",x"8e"),
  1768 => (x"c0",x"48",x"f0",x"fe"),
  1769 => (x"79",x"09",x"cd",x"78"),
  1770 => (x"1e",x"4f",x"26",x"09"),
  1771 => (x"49",x"d4",x"ee",x"c1"),
  1772 => (x"4f",x"26",x"87",x"ed"),
  1773 => (x"bf",x"f0",x"fe",x"1e"),
  1774 => (x"1e",x"4f",x"26",x"48"),
  1775 => (x"c1",x"48",x"f0",x"fe"),
  1776 => (x"1e",x"4f",x"26",x"78"),
  1777 => (x"c0",x"48",x"f0",x"fe"),
  1778 => (x"1e",x"4f",x"26",x"78"),
  1779 => (x"52",x"c0",x"4a",x"71"),
  1780 => (x"0e",x"4f",x"26",x"51"),
  1781 => (x"5d",x"5c",x"5b",x"5e"),
  1782 => (x"71",x"86",x"f4",x"0e"),
  1783 => (x"7e",x"6d",x"97",x"4d"),
  1784 => (x"97",x"4c",x"a5",x"c1"),
  1785 => (x"a6",x"c8",x"48",x"6c"),
  1786 => (x"c4",x"48",x"6e",x"58"),
  1787 => (x"c5",x"05",x"a8",x"66"),
  1788 => (x"c0",x"48",x"ff",x"87"),
  1789 => (x"ca",x"ff",x"87",x"e6"),
  1790 => (x"49",x"a5",x"c2",x"87"),
  1791 => (x"71",x"4b",x"6c",x"97"),
  1792 => (x"6b",x"97",x"4b",x"a3"),
  1793 => (x"7e",x"6c",x"97",x"4b"),
  1794 => (x"80",x"c1",x"48",x"6e"),
  1795 => (x"c7",x"58",x"a6",x"c8"),
  1796 => (x"58",x"a6",x"cc",x"98"),
  1797 => (x"fe",x"7c",x"97",x"70"),
  1798 => (x"48",x"73",x"87",x"e1"),
  1799 => (x"4d",x"26",x"8e",x"f4"),
  1800 => (x"4b",x"26",x"4c",x"26"),
  1801 => (x"5e",x"0e",x"4f",x"26"),
  1802 => (x"f4",x"0e",x"5c",x"5b"),
  1803 => (x"d8",x"4c",x"71",x"86"),
  1804 => (x"ff",x"c3",x"4a",x"66"),
  1805 => (x"4b",x"a4",x"c2",x"9a"),
  1806 => (x"73",x"49",x"6c",x"97"),
  1807 => (x"51",x"72",x"49",x"a1"),
  1808 => (x"6e",x"7e",x"6c",x"97"),
  1809 => (x"c8",x"80",x"c1",x"48"),
  1810 => (x"98",x"c7",x"58",x"a6"),
  1811 => (x"70",x"58",x"a6",x"cc"),
  1812 => (x"26",x"8e",x"f4",x"54"),
  1813 => (x"26",x"4b",x"26",x"4c"),
  1814 => (x"86",x"fc",x"1e",x"4f"),
  1815 => (x"e0",x"87",x"e4",x"fd"),
  1816 => (x"c0",x"49",x"4a",x"bf"),
  1817 => (x"02",x"99",x"c0",x"e0"),
  1818 => (x"1e",x"72",x"87",x"cb"),
  1819 => (x"49",x"f4",x"f4",x"c2"),
  1820 => (x"c4",x"87",x"f3",x"fe"),
  1821 => (x"87",x"fc",x"fc",x"86"),
  1822 => (x"fe",x"fc",x"7e",x"70"),
  1823 => (x"26",x"8e",x"fc",x"87"),
  1824 => (x"f4",x"c2",x"1e",x"4f"),
  1825 => (x"c2",x"fd",x"49",x"f4"),
  1826 => (x"d9",x"f1",x"c1",x"87"),
  1827 => (x"87",x"cf",x"fc",x"49"),
  1828 => (x"26",x"87",x"ed",x"c3"),
  1829 => (x"5b",x"5e",x"0e",x"4f"),
  1830 => (x"fc",x"0e",x"5d",x"5c"),
  1831 => (x"ff",x"7e",x"71",x"86"),
  1832 => (x"f4",x"c2",x"4d",x"d4"),
  1833 => (x"ea",x"fc",x"49",x"f4"),
  1834 => (x"c0",x"4b",x"70",x"87"),
  1835 => (x"c2",x"04",x"ab",x"b7"),
  1836 => (x"f0",x"c3",x"87",x"f8"),
  1837 => (x"87",x"c9",x"05",x"ab"),
  1838 => (x"48",x"f8",x"f5",x"c1"),
  1839 => (x"d9",x"c2",x"78",x"c1"),
  1840 => (x"ab",x"e0",x"c3",x"87"),
  1841 => (x"c1",x"87",x"c9",x"05"),
  1842 => (x"c1",x"48",x"fc",x"f5"),
  1843 => (x"87",x"ca",x"c2",x"78"),
  1844 => (x"bf",x"fc",x"f5",x"c1"),
  1845 => (x"c2",x"87",x"c6",x"02"),
  1846 => (x"c2",x"4c",x"a3",x"c0"),
  1847 => (x"c1",x"4c",x"73",x"87"),
  1848 => (x"02",x"bf",x"f8",x"f5"),
  1849 => (x"74",x"87",x"e0",x"c0"),
  1850 => (x"29",x"b7",x"c4",x"49"),
  1851 => (x"d4",x"f7",x"c1",x"91"),
  1852 => (x"cf",x"4a",x"74",x"81"),
  1853 => (x"c1",x"92",x"c2",x"9a"),
  1854 => (x"70",x"30",x"72",x"48"),
  1855 => (x"72",x"ba",x"ff",x"4a"),
  1856 => (x"70",x"98",x"69",x"48"),
  1857 => (x"74",x"87",x"db",x"79"),
  1858 => (x"29",x"b7",x"c4",x"49"),
  1859 => (x"d4",x"f7",x"c1",x"91"),
  1860 => (x"cf",x"4a",x"74",x"81"),
  1861 => (x"c3",x"92",x"c2",x"9a"),
  1862 => (x"70",x"30",x"72",x"48"),
  1863 => (x"b0",x"69",x"48",x"4a"),
  1864 => (x"05",x"6e",x"79",x"70"),
  1865 => (x"ff",x"87",x"e7",x"c0"),
  1866 => (x"e1",x"c8",x"48",x"d0"),
  1867 => (x"c1",x"7d",x"c5",x"78"),
  1868 => (x"02",x"bf",x"fc",x"f5"),
  1869 => (x"e0",x"c3",x"87",x"c3"),
  1870 => (x"f8",x"f5",x"c1",x"7d"),
  1871 => (x"87",x"c3",x"02",x"bf"),
  1872 => (x"73",x"7d",x"f0",x"c3"),
  1873 => (x"48",x"d0",x"ff",x"7d"),
  1874 => (x"c0",x"78",x"e1",x"c8"),
  1875 => (x"f5",x"c1",x"78",x"e0"),
  1876 => (x"78",x"c0",x"48",x"fc"),
  1877 => (x"48",x"f8",x"f5",x"c1"),
  1878 => (x"f4",x"c2",x"78",x"c0"),
  1879 => (x"f2",x"f9",x"49",x"f4"),
  1880 => (x"c0",x"4b",x"70",x"87"),
  1881 => (x"fd",x"03",x"ab",x"b7"),
  1882 => (x"48",x"c0",x"87",x"c8"),
  1883 => (x"4d",x"26",x"8e",x"fc"),
  1884 => (x"4b",x"26",x"4c",x"26"),
  1885 => (x"00",x"00",x"4f",x"26"),
  1886 => (x"00",x"00",x"00",x"00"),
  1887 => (x"00",x"00",x"00",x"00"),
  1888 => (x"72",x"4a",x"c0",x"1e"),
  1889 => (x"c1",x"91",x"c4",x"49"),
  1890 => (x"c0",x"81",x"d4",x"f7"),
  1891 => (x"d0",x"82",x"c1",x"79"),
  1892 => (x"ee",x"04",x"aa",x"b7"),
  1893 => (x"0e",x"4f",x"26",x"87"),
  1894 => (x"5d",x"5c",x"5b",x"5e"),
  1895 => (x"f8",x"4d",x"71",x"0e"),
  1896 => (x"4a",x"75",x"87",x"e1"),
  1897 => (x"92",x"2a",x"b7",x"c4"),
  1898 => (x"82",x"d4",x"f7",x"c1"),
  1899 => (x"9c",x"cf",x"4c",x"75"),
  1900 => (x"49",x"6a",x"94",x"c2"),
  1901 => (x"c3",x"2b",x"74",x"4b"),
  1902 => (x"74",x"48",x"c2",x"9b"),
  1903 => (x"ff",x"4c",x"70",x"30"),
  1904 => (x"71",x"48",x"74",x"bc"),
  1905 => (x"f7",x"7a",x"70",x"98"),
  1906 => (x"48",x"73",x"87",x"f1"),
  1907 => (x"4c",x"26",x"4d",x"26"),
  1908 => (x"4f",x"26",x"4b",x"26"),
  1909 => (x"00",x"00",x"00",x"00"),
  1910 => (x"00",x"00",x"00",x"00"),
  1911 => (x"00",x"00",x"00",x"00"),
  1912 => (x"00",x"00",x"00",x"00"),
  1913 => (x"00",x"00",x"00",x"00"),
  1914 => (x"00",x"00",x"00",x"00"),
  1915 => (x"00",x"00",x"00",x"00"),
  1916 => (x"00",x"00",x"00",x"00"),
  1917 => (x"00",x"00",x"00",x"00"),
  1918 => (x"00",x"00",x"00",x"00"),
  1919 => (x"00",x"00",x"00",x"00"),
  1920 => (x"00",x"00",x"00",x"00"),
  1921 => (x"00",x"00",x"00",x"00"),
  1922 => (x"00",x"00",x"00",x"00"),
  1923 => (x"00",x"00",x"00",x"00"),
  1924 => (x"00",x"00",x"00",x"00"),
  1925 => (x"48",x"d0",x"ff",x"1e"),
  1926 => (x"71",x"78",x"e1",x"c8"),
  1927 => (x"08",x"d4",x"ff",x"48"),
  1928 => (x"1e",x"4f",x"26",x"78"),
  1929 => (x"c8",x"48",x"d0",x"ff"),
  1930 => (x"48",x"71",x"78",x"e1"),
  1931 => (x"78",x"08",x"d4",x"ff"),
  1932 => (x"ff",x"48",x"66",x"c4"),
  1933 => (x"26",x"78",x"08",x"d4"),
  1934 => (x"4a",x"71",x"1e",x"4f"),
  1935 => (x"1e",x"49",x"66",x"c4"),
  1936 => (x"de",x"ff",x"49",x"72"),
  1937 => (x"48",x"d0",x"ff",x"87"),
  1938 => (x"fc",x"78",x"e0",x"c0"),
  1939 => (x"1e",x"4f",x"26",x"8e"),
  1940 => (x"4b",x"71",x"1e",x"73"),
  1941 => (x"1e",x"49",x"66",x"c8"),
  1942 => (x"e0",x"c1",x"4a",x"73"),
  1943 => (x"d8",x"ff",x"49",x"a2"),
  1944 => (x"26",x"8e",x"fc",x"87"),
  1945 => (x"1e",x"4f",x"26",x"4b"),
  1946 => (x"c8",x"48",x"d0",x"ff"),
  1947 => (x"48",x"71",x"78",x"c9"),
  1948 => (x"78",x"08",x"d4",x"ff"),
  1949 => (x"71",x"1e",x"4f",x"26"),
  1950 => (x"87",x"eb",x"49",x"4a"),
  1951 => (x"c8",x"48",x"d0",x"ff"),
  1952 => (x"1e",x"4f",x"26",x"78"),
  1953 => (x"4b",x"71",x"1e",x"73"),
  1954 => (x"bf",x"cc",x"f5",x"c2"),
  1955 => (x"c2",x"87",x"c3",x"02"),
  1956 => (x"d0",x"ff",x"87",x"eb"),
  1957 => (x"78",x"c9",x"c8",x"48"),
  1958 => (x"e0",x"c0",x"48",x"73"),
  1959 => (x"08",x"d4",x"ff",x"b0"),
  1960 => (x"c0",x"f5",x"c2",x"78"),
  1961 => (x"c8",x"78",x"c0",x"48"),
  1962 => (x"87",x"c5",x"02",x"66"),
  1963 => (x"c2",x"49",x"ff",x"c3"),
  1964 => (x"c2",x"49",x"c0",x"87"),
  1965 => (x"cc",x"59",x"c8",x"f5"),
  1966 => (x"87",x"c6",x"02",x"66"),
  1967 => (x"4a",x"d5",x"d5",x"c5"),
  1968 => (x"ff",x"cf",x"87",x"c4"),
  1969 => (x"f5",x"c2",x"4a",x"ff"),
  1970 => (x"f5",x"c2",x"5a",x"cc"),
  1971 => (x"78",x"c1",x"48",x"cc"),
  1972 => (x"4f",x"26",x"4b",x"26"),
  1973 => (x"5c",x"5b",x"5e",x"0e"),
  1974 => (x"4d",x"71",x"0e",x"5d"),
  1975 => (x"bf",x"c8",x"f5",x"c2"),
  1976 => (x"02",x"9d",x"75",x"4b"),
  1977 => (x"c8",x"49",x"87",x"cb"),
  1978 => (x"fc",x"f9",x"c1",x"91"),
  1979 => (x"c4",x"82",x"71",x"4a"),
  1980 => (x"fc",x"fd",x"c1",x"87"),
  1981 => (x"12",x"4c",x"c0",x"4a"),
  1982 => (x"c2",x"99",x"73",x"49"),
  1983 => (x"48",x"bf",x"c4",x"f5"),
  1984 => (x"d4",x"ff",x"b8",x"71"),
  1985 => (x"b7",x"c1",x"78",x"08"),
  1986 => (x"b7",x"c8",x"84",x"2b"),
  1987 => (x"87",x"e7",x"04",x"ac"),
  1988 => (x"bf",x"c0",x"f5",x"c2"),
  1989 => (x"c2",x"80",x"c8",x"48"),
  1990 => (x"26",x"58",x"c4",x"f5"),
  1991 => (x"26",x"4c",x"26",x"4d"),
  1992 => (x"1e",x"4f",x"26",x"4b"),
  1993 => (x"4b",x"71",x"1e",x"73"),
  1994 => (x"02",x"9a",x"4a",x"13"),
  1995 => (x"49",x"72",x"87",x"cb"),
  1996 => (x"13",x"87",x"e1",x"fe"),
  1997 => (x"f5",x"05",x"9a",x"4a"),
  1998 => (x"26",x"4b",x"26",x"87"),
  1999 => (x"f5",x"c2",x"1e",x"4f"),
  2000 => (x"c2",x"49",x"bf",x"c0"),
  2001 => (x"c1",x"48",x"c0",x"f5"),
  2002 => (x"c0",x"c4",x"78",x"a1"),
  2003 => (x"db",x"03",x"a9",x"b7"),
  2004 => (x"48",x"d4",x"ff",x"87"),
  2005 => (x"bf",x"c4",x"f5",x"c2"),
  2006 => (x"c0",x"f5",x"c2",x"78"),
  2007 => (x"f5",x"c2",x"49",x"bf"),
  2008 => (x"a1",x"c1",x"48",x"c0"),
  2009 => (x"b7",x"c0",x"c4",x"78"),
  2010 => (x"87",x"e5",x"04",x"a9"),
  2011 => (x"c8",x"48",x"d0",x"ff"),
  2012 => (x"cc",x"f5",x"c2",x"78"),
  2013 => (x"26",x"78",x"c0",x"48"),
  2014 => (x"00",x"00",x"00",x"4f"),
  2015 => (x"00",x"00",x"00",x"00"),
  2016 => (x"00",x"00",x"00",x"00"),
  2017 => (x"5f",x"00",x"00",x"00"),
  2018 => (x"00",x"00",x"00",x"5f"),
  2019 => (x"00",x"03",x"03",x"00"),
  2020 => (x"00",x"00",x"03",x"03"),
  2021 => (x"14",x"7f",x"7f",x"14"),
  2022 => (x"00",x"14",x"7f",x"7f"),
  2023 => (x"6b",x"2e",x"24",x"00"),
  2024 => (x"00",x"12",x"3a",x"6b"),
  2025 => (x"18",x"36",x"6a",x"4c"),
  2026 => (x"00",x"32",x"56",x"6c"),
  2027 => (x"59",x"4f",x"7e",x"30"),
  2028 => (x"40",x"68",x"3a",x"77"),
  2029 => (x"07",x"04",x"00",x"00"),
  2030 => (x"00",x"00",x"00",x"03"),
  2031 => (x"3e",x"1c",x"00",x"00"),
  2032 => (x"00",x"00",x"41",x"63"),
  2033 => (x"63",x"41",x"00",x"00"),
  2034 => (x"00",x"00",x"1c",x"3e"),
  2035 => (x"1c",x"3e",x"2a",x"08"),
  2036 => (x"08",x"2a",x"3e",x"1c"),
  2037 => (x"3e",x"08",x"08",x"00"),
  2038 => (x"00",x"08",x"08",x"3e"),
  2039 => (x"e0",x"80",x"00",x"00"),
  2040 => (x"00",x"00",x"00",x"60"),
  2041 => (x"08",x"08",x"08",x"00"),
  2042 => (x"00",x"08",x"08",x"08"),
  2043 => (x"60",x"00",x"00",x"00"),
  2044 => (x"00",x"00",x"00",x"60"),
  2045 => (x"18",x"30",x"60",x"40"),
  2046 => (x"01",x"03",x"06",x"0c"),
  2047 => (x"59",x"7f",x"3e",x"00"),
  2048 => (x"00",x"3e",x"7f",x"4d"),
  2049 => (x"7f",x"06",x"04",x"00"),
  2050 => (x"00",x"00",x"00",x"7f"),
  2051 => (x"71",x"63",x"42",x"00"),
  2052 => (x"00",x"46",x"4f",x"59"),
  2053 => (x"49",x"63",x"22",x"00"),
  2054 => (x"00",x"36",x"7f",x"49"),
  2055 => (x"13",x"16",x"1c",x"18"),
  2056 => (x"00",x"10",x"7f",x"7f"),
  2057 => (x"45",x"67",x"27",x"00"),
  2058 => (x"00",x"39",x"7d",x"45"),
  2059 => (x"4b",x"7e",x"3c",x"00"),
  2060 => (x"00",x"30",x"79",x"49"),
  2061 => (x"71",x"01",x"01",x"00"),
  2062 => (x"00",x"07",x"0f",x"79"),
  2063 => (x"49",x"7f",x"36",x"00"),
  2064 => (x"00",x"36",x"7f",x"49"),
  2065 => (x"49",x"4f",x"06",x"00"),
  2066 => (x"00",x"1e",x"3f",x"69"),
  2067 => (x"66",x"00",x"00",x"00"),
  2068 => (x"00",x"00",x"00",x"66"),
  2069 => (x"e6",x"80",x"00",x"00"),
  2070 => (x"00",x"00",x"00",x"66"),
  2071 => (x"14",x"08",x"08",x"00"),
  2072 => (x"00",x"22",x"22",x"14"),
  2073 => (x"14",x"14",x"14",x"00"),
  2074 => (x"00",x"14",x"14",x"14"),
  2075 => (x"14",x"22",x"22",x"00"),
  2076 => (x"00",x"08",x"08",x"14"),
  2077 => (x"51",x"03",x"02",x"00"),
  2078 => (x"00",x"06",x"0f",x"59"),
  2079 => (x"5d",x"41",x"7f",x"3e"),
  2080 => (x"00",x"1e",x"1f",x"55"),
  2081 => (x"09",x"7f",x"7e",x"00"),
  2082 => (x"00",x"7e",x"7f",x"09"),
  2083 => (x"49",x"7f",x"7f",x"00"),
  2084 => (x"00",x"36",x"7f",x"49"),
  2085 => (x"63",x"3e",x"1c",x"00"),
  2086 => (x"00",x"41",x"41",x"41"),
  2087 => (x"41",x"7f",x"7f",x"00"),
  2088 => (x"00",x"1c",x"3e",x"63"),
  2089 => (x"49",x"7f",x"7f",x"00"),
  2090 => (x"00",x"41",x"41",x"49"),
  2091 => (x"09",x"7f",x"7f",x"00"),
  2092 => (x"00",x"01",x"01",x"09"),
  2093 => (x"41",x"7f",x"3e",x"00"),
  2094 => (x"00",x"7a",x"7b",x"49"),
  2095 => (x"08",x"7f",x"7f",x"00"),
  2096 => (x"00",x"7f",x"7f",x"08"),
  2097 => (x"7f",x"41",x"00",x"00"),
  2098 => (x"00",x"00",x"41",x"7f"),
  2099 => (x"40",x"60",x"20",x"00"),
  2100 => (x"00",x"3f",x"7f",x"40"),
  2101 => (x"1c",x"08",x"7f",x"7f"),
  2102 => (x"00",x"41",x"63",x"36"),
  2103 => (x"40",x"7f",x"7f",x"00"),
  2104 => (x"00",x"40",x"40",x"40"),
  2105 => (x"0c",x"06",x"7f",x"7f"),
  2106 => (x"00",x"7f",x"7f",x"06"),
  2107 => (x"0c",x"06",x"7f",x"7f"),
  2108 => (x"00",x"7f",x"7f",x"18"),
  2109 => (x"41",x"7f",x"3e",x"00"),
  2110 => (x"00",x"3e",x"7f",x"41"),
  2111 => (x"09",x"7f",x"7f",x"00"),
  2112 => (x"00",x"06",x"0f",x"09"),
  2113 => (x"61",x"41",x"7f",x"3e"),
  2114 => (x"00",x"40",x"7e",x"7f"),
  2115 => (x"09",x"7f",x"7f",x"00"),
  2116 => (x"00",x"66",x"7f",x"19"),
  2117 => (x"4d",x"6f",x"26",x"00"),
  2118 => (x"00",x"32",x"7b",x"59"),
  2119 => (x"7f",x"01",x"01",x"00"),
  2120 => (x"00",x"01",x"01",x"7f"),
  2121 => (x"40",x"7f",x"3f",x"00"),
  2122 => (x"00",x"3f",x"7f",x"40"),
  2123 => (x"70",x"3f",x"0f",x"00"),
  2124 => (x"00",x"0f",x"3f",x"70"),
  2125 => (x"18",x"30",x"7f",x"7f"),
  2126 => (x"00",x"7f",x"7f",x"30"),
  2127 => (x"1c",x"36",x"63",x"41"),
  2128 => (x"41",x"63",x"36",x"1c"),
  2129 => (x"7c",x"06",x"03",x"01"),
  2130 => (x"01",x"03",x"06",x"7c"),
  2131 => (x"4d",x"59",x"71",x"61"),
  2132 => (x"00",x"41",x"43",x"47"),
  2133 => (x"7f",x"7f",x"00",x"00"),
  2134 => (x"00",x"00",x"41",x"41"),
  2135 => (x"0c",x"06",x"03",x"01"),
  2136 => (x"40",x"60",x"30",x"18"),
  2137 => (x"41",x"41",x"00",x"00"),
  2138 => (x"00",x"00",x"7f",x"7f"),
  2139 => (x"03",x"06",x"0c",x"08"),
  2140 => (x"00",x"08",x"0c",x"06"),
  2141 => (x"80",x"80",x"80",x"80"),
  2142 => (x"00",x"80",x"80",x"80"),
  2143 => (x"03",x"00",x"00",x"00"),
  2144 => (x"00",x"00",x"04",x"07"),
  2145 => (x"54",x"74",x"20",x"00"),
  2146 => (x"00",x"78",x"7c",x"54"),
  2147 => (x"44",x"7f",x"7f",x"00"),
  2148 => (x"00",x"38",x"7c",x"44"),
  2149 => (x"44",x"7c",x"38",x"00"),
  2150 => (x"00",x"00",x"44",x"44"),
  2151 => (x"44",x"7c",x"38",x"00"),
  2152 => (x"00",x"7f",x"7f",x"44"),
  2153 => (x"54",x"7c",x"38",x"00"),
  2154 => (x"00",x"18",x"5c",x"54"),
  2155 => (x"7f",x"7e",x"04",x"00"),
  2156 => (x"00",x"00",x"05",x"05"),
  2157 => (x"a4",x"bc",x"18",x"00"),
  2158 => (x"00",x"7c",x"fc",x"a4"),
  2159 => (x"04",x"7f",x"7f",x"00"),
  2160 => (x"00",x"78",x"7c",x"04"),
  2161 => (x"3d",x"00",x"00",x"00"),
  2162 => (x"00",x"00",x"40",x"7d"),
  2163 => (x"80",x"80",x"80",x"00"),
  2164 => (x"00",x"00",x"7d",x"fd"),
  2165 => (x"10",x"7f",x"7f",x"00"),
  2166 => (x"00",x"44",x"6c",x"38"),
  2167 => (x"3f",x"00",x"00",x"00"),
  2168 => (x"00",x"00",x"40",x"7f"),
  2169 => (x"18",x"0c",x"7c",x"7c"),
  2170 => (x"00",x"78",x"7c",x"0c"),
  2171 => (x"04",x"7c",x"7c",x"00"),
  2172 => (x"00",x"78",x"7c",x"04"),
  2173 => (x"44",x"7c",x"38",x"00"),
  2174 => (x"00",x"38",x"7c",x"44"),
  2175 => (x"24",x"fc",x"fc",x"00"),
  2176 => (x"00",x"18",x"3c",x"24"),
  2177 => (x"24",x"3c",x"18",x"00"),
  2178 => (x"00",x"fc",x"fc",x"24"),
  2179 => (x"04",x"7c",x"7c",x"00"),
  2180 => (x"00",x"08",x"0c",x"04"),
  2181 => (x"54",x"5c",x"48",x"00"),
  2182 => (x"00",x"20",x"74",x"54"),
  2183 => (x"7f",x"3f",x"04",x"00"),
  2184 => (x"00",x"00",x"44",x"44"),
  2185 => (x"40",x"7c",x"3c",x"00"),
  2186 => (x"00",x"7c",x"7c",x"40"),
  2187 => (x"60",x"3c",x"1c",x"00"),
  2188 => (x"00",x"1c",x"3c",x"60"),
  2189 => (x"30",x"60",x"7c",x"3c"),
  2190 => (x"00",x"3c",x"7c",x"60"),
  2191 => (x"10",x"38",x"6c",x"44"),
  2192 => (x"00",x"44",x"6c",x"38"),
  2193 => (x"e0",x"bc",x"1c",x"00"),
  2194 => (x"00",x"1c",x"3c",x"60"),
  2195 => (x"74",x"64",x"44",x"00"),
  2196 => (x"00",x"44",x"4c",x"5c"),
  2197 => (x"3e",x"08",x"08",x"00"),
  2198 => (x"00",x"41",x"41",x"77"),
  2199 => (x"7f",x"00",x"00",x"00"),
  2200 => (x"00",x"00",x"00",x"7f"),
  2201 => (x"77",x"41",x"41",x"00"),
  2202 => (x"00",x"08",x"08",x"3e"),
  2203 => (x"03",x"01",x"01",x"02"),
  2204 => (x"00",x"01",x"02",x"02"),
  2205 => (x"7f",x"7f",x"7f",x"7f"),
  2206 => (x"00",x"7f",x"7f",x"7f"),
  2207 => (x"1c",x"1c",x"08",x"08"),
  2208 => (x"7f",x"7f",x"3e",x"3e"),
  2209 => (x"3e",x"3e",x"7f",x"7f"),
  2210 => (x"08",x"08",x"1c",x"1c"),
  2211 => (x"7c",x"18",x"10",x"00"),
  2212 => (x"00",x"10",x"18",x"7c"),
  2213 => (x"7c",x"30",x"10",x"00"),
  2214 => (x"00",x"10",x"30",x"7c"),
  2215 => (x"60",x"60",x"30",x"10"),
  2216 => (x"00",x"06",x"1e",x"78"),
  2217 => (x"18",x"3c",x"66",x"42"),
  2218 => (x"00",x"42",x"66",x"3c"),
  2219 => (x"c2",x"6a",x"38",x"78"),
  2220 => (x"00",x"38",x"6c",x"c6"),
  2221 => (x"60",x"00",x"00",x"60"),
  2222 => (x"00",x"60",x"00",x"00"),
  2223 => (x"5c",x"5b",x"5e",x"0e"),
  2224 => (x"86",x"fc",x"0e",x"5d"),
  2225 => (x"f5",x"c2",x"7e",x"71"),
  2226 => (x"c0",x"4c",x"bf",x"d4"),
  2227 => (x"c4",x"1e",x"c0",x"4b"),
  2228 => (x"c4",x"02",x"ab",x"66"),
  2229 => (x"c2",x"4d",x"c0",x"87"),
  2230 => (x"75",x"4d",x"c1",x"87"),
  2231 => (x"ee",x"49",x"73",x"1e"),
  2232 => (x"86",x"c8",x"87",x"e1"),
  2233 => (x"ef",x"49",x"e0",x"c0"),
  2234 => (x"a4",x"c4",x"87",x"ea"),
  2235 => (x"f0",x"49",x"6a",x"4a"),
  2236 => (x"c8",x"f1",x"87",x"f1"),
  2237 => (x"c1",x"84",x"cc",x"87"),
  2238 => (x"ab",x"b7",x"c8",x"83"),
  2239 => (x"87",x"cd",x"ff",x"04"),
  2240 => (x"4d",x"26",x"8e",x"fc"),
  2241 => (x"4b",x"26",x"4c",x"26"),
  2242 => (x"71",x"1e",x"4f",x"26"),
  2243 => (x"d8",x"f5",x"c2",x"4a"),
  2244 => (x"d8",x"f5",x"c2",x"5a"),
  2245 => (x"49",x"78",x"c7",x"48"),
  2246 => (x"26",x"87",x"e1",x"fe"),
  2247 => (x"1e",x"73",x"1e",x"4f"),
  2248 => (x"b7",x"c0",x"4a",x"71"),
  2249 => (x"87",x"d3",x"03",x"aa"),
  2250 => (x"bf",x"f8",x"d9",x"c2"),
  2251 => (x"c1",x"87",x"c4",x"05"),
  2252 => (x"c0",x"87",x"c2",x"4b"),
  2253 => (x"fc",x"d9",x"c2",x"4b"),
  2254 => (x"c2",x"87",x"c4",x"5b"),
  2255 => (x"fc",x"5a",x"fc",x"d9"),
  2256 => (x"f8",x"d9",x"c2",x"48"),
  2257 => (x"c1",x"4a",x"78",x"bf"),
  2258 => (x"a2",x"c0",x"c1",x"9a"),
  2259 => (x"87",x"e6",x"ec",x"49"),
  2260 => (x"4f",x"26",x"4b",x"26"),
  2261 => (x"c4",x"4a",x"71",x"1e"),
  2262 => (x"49",x"72",x"1e",x"66"),
  2263 => (x"fc",x"87",x"f0",x"eb"),
  2264 => (x"1e",x"4f",x"26",x"8e"),
  2265 => (x"c3",x"48",x"d4",x"ff"),
  2266 => (x"d0",x"ff",x"78",x"ff"),
  2267 => (x"78",x"e1",x"c0",x"48"),
  2268 => (x"c1",x"48",x"d4",x"ff"),
  2269 => (x"c4",x"48",x"71",x"78"),
  2270 => (x"08",x"d4",x"ff",x"30"),
  2271 => (x"48",x"d0",x"ff",x"78"),
  2272 => (x"26",x"78",x"e0",x"c0"),
  2273 => (x"5b",x"5e",x"0e",x"4f"),
  2274 => (x"ec",x"0e",x"5d",x"5c"),
  2275 => (x"48",x"a6",x"c8",x"86"),
  2276 => (x"c4",x"7e",x"78",x"c0"),
  2277 => (x"78",x"bf",x"ec",x"80"),
  2278 => (x"f5",x"c2",x"80",x"f8"),
  2279 => (x"e8",x"78",x"bf",x"d4"),
  2280 => (x"d9",x"c2",x"4c",x"bf"),
  2281 => (x"e3",x"49",x"bf",x"f8"),
  2282 => (x"ee",x"cb",x"87",x"eb"),
  2283 => (x"87",x"cc",x"cb",x"49"),
  2284 => (x"c7",x"58",x"a6",x"d4"),
  2285 => (x"87",x"df",x"e7",x"49"),
  2286 => (x"c9",x"05",x"98",x"70"),
  2287 => (x"49",x"66",x"cc",x"87"),
  2288 => (x"c1",x"02",x"99",x"c1"),
  2289 => (x"66",x"d0",x"87",x"c4"),
  2290 => (x"ec",x"7e",x"c1",x"4d"),
  2291 => (x"d9",x"c2",x"4b",x"bf"),
  2292 => (x"e2",x"49",x"bf",x"f8"),
  2293 => (x"49",x"75",x"87",x"ff"),
  2294 => (x"70",x"87",x"ed",x"ca"),
  2295 => (x"87",x"d7",x"02",x"98"),
  2296 => (x"bf",x"e0",x"d9",x"c2"),
  2297 => (x"c2",x"b9",x"c1",x"49"),
  2298 => (x"71",x"59",x"e4",x"d9"),
  2299 => (x"cb",x"87",x"f4",x"fd"),
  2300 => (x"c7",x"ca",x"49",x"ee"),
  2301 => (x"c7",x"4d",x"70",x"87"),
  2302 => (x"87",x"db",x"e6",x"49"),
  2303 => (x"ff",x"05",x"98",x"70"),
  2304 => (x"49",x"73",x"87",x"c7"),
  2305 => (x"fe",x"05",x"99",x"c1"),
  2306 => (x"02",x"6e",x"87",x"ff"),
  2307 => (x"c2",x"87",x"e3",x"c0"),
  2308 => (x"4a",x"bf",x"f8",x"d9"),
  2309 => (x"d9",x"c2",x"ba",x"c1"),
  2310 => (x"0a",x"fc",x"5a",x"fc"),
  2311 => (x"9a",x"c1",x"0a",x"7a"),
  2312 => (x"49",x"a2",x"c0",x"c1"),
  2313 => (x"c1",x"87",x"cf",x"e9"),
  2314 => (x"ea",x"e5",x"49",x"da"),
  2315 => (x"48",x"a6",x"c8",x"87"),
  2316 => (x"d9",x"c2",x"78",x"c1"),
  2317 => (x"c1",x"05",x"bf",x"f8"),
  2318 => (x"c0",x"c8",x"87",x"c5"),
  2319 => (x"d9",x"c2",x"4d",x"c0"),
  2320 => (x"49",x"13",x"4b",x"e4"),
  2321 => (x"87",x"cf",x"e5",x"49"),
  2322 => (x"c2",x"02",x"98",x"70"),
  2323 => (x"c1",x"b4",x"75",x"87"),
  2324 => (x"ff",x"05",x"2d",x"b7"),
  2325 => (x"49",x"74",x"87",x"ec"),
  2326 => (x"71",x"99",x"ff",x"c3"),
  2327 => (x"fb",x"49",x"c0",x"1e"),
  2328 => (x"49",x"74",x"87",x"f2"),
  2329 => (x"71",x"29",x"b7",x"c8"),
  2330 => (x"fb",x"49",x"c1",x"1e"),
  2331 => (x"86",x"c8",x"87",x"e6"),
  2332 => (x"e4",x"49",x"fd",x"c3"),
  2333 => (x"fa",x"c3",x"87",x"e1"),
  2334 => (x"87",x"db",x"e4",x"49"),
  2335 => (x"74",x"87",x"d4",x"c7"),
  2336 => (x"99",x"ff",x"c3",x"49"),
  2337 => (x"71",x"2c",x"b7",x"c8"),
  2338 => (x"02",x"9c",x"74",x"b4"),
  2339 => (x"d9",x"c2",x"87",x"df"),
  2340 => (x"c7",x"49",x"bf",x"f4"),
  2341 => (x"98",x"70",x"87",x"f2"),
  2342 => (x"87",x"c4",x"c0",x"05"),
  2343 => (x"87",x"d3",x"4c",x"c0"),
  2344 => (x"c7",x"49",x"e0",x"c2"),
  2345 => (x"d9",x"c2",x"87",x"d6"),
  2346 => (x"c6",x"c0",x"58",x"f8"),
  2347 => (x"f4",x"d9",x"c2",x"87"),
  2348 => (x"74",x"78",x"c0",x"48"),
  2349 => (x"05",x"99",x"c8",x"49"),
  2350 => (x"c3",x"87",x"ce",x"c0"),
  2351 => (x"d6",x"e3",x"49",x"f5"),
  2352 => (x"c2",x"49",x"70",x"87"),
  2353 => (x"e7",x"c0",x"02",x"99"),
  2354 => (x"d8",x"f5",x"c2",x"87"),
  2355 => (x"ca",x"c0",x"02",x"bf"),
  2356 => (x"88",x"c1",x"48",x"87"),
  2357 => (x"58",x"dc",x"f5",x"c2"),
  2358 => (x"c4",x"87",x"d0",x"c0"),
  2359 => (x"e0",x"c1",x"4a",x"66"),
  2360 => (x"c0",x"02",x"6a",x"82"),
  2361 => (x"ff",x"4b",x"87",x"c5"),
  2362 => (x"c8",x"0f",x"73",x"49"),
  2363 => (x"78",x"c1",x"48",x"a6"),
  2364 => (x"99",x"c4",x"49",x"74"),
  2365 => (x"87",x"ce",x"c0",x"05"),
  2366 => (x"e2",x"49",x"f2",x"c3"),
  2367 => (x"49",x"70",x"87",x"d9"),
  2368 => (x"c0",x"02",x"99",x"c2"),
  2369 => (x"f5",x"c2",x"87",x"f0"),
  2370 => (x"48",x"7e",x"bf",x"d8"),
  2371 => (x"03",x"a8",x"b7",x"c7"),
  2372 => (x"6e",x"87",x"cb",x"c0"),
  2373 => (x"c2",x"80",x"c1",x"48"),
  2374 => (x"c0",x"58",x"dc",x"f5"),
  2375 => (x"66",x"c4",x"87",x"d3"),
  2376 => (x"80",x"e0",x"c1",x"48"),
  2377 => (x"bf",x"6e",x"7e",x"70"),
  2378 => (x"87",x"c5",x"c0",x"02"),
  2379 => (x"73",x"49",x"fe",x"4b"),
  2380 => (x"48",x"a6",x"c8",x"0f"),
  2381 => (x"fd",x"c3",x"78",x"c1"),
  2382 => (x"87",x"db",x"e1",x"49"),
  2383 => (x"99",x"c2",x"49",x"70"),
  2384 => (x"87",x"e9",x"c0",x"02"),
  2385 => (x"bf",x"d8",x"f5",x"c2"),
  2386 => (x"87",x"c9",x"c0",x"02"),
  2387 => (x"48",x"d8",x"f5",x"c2"),
  2388 => (x"d3",x"c0",x"78",x"c0"),
  2389 => (x"48",x"66",x"c4",x"87"),
  2390 => (x"70",x"80",x"e0",x"c1"),
  2391 => (x"02",x"bf",x"6e",x"7e"),
  2392 => (x"4b",x"87",x"c5",x"c0"),
  2393 => (x"0f",x"73",x"49",x"fd"),
  2394 => (x"c1",x"48",x"a6",x"c8"),
  2395 => (x"49",x"fa",x"c3",x"78"),
  2396 => (x"70",x"87",x"e4",x"e0"),
  2397 => (x"02",x"99",x"c2",x"49"),
  2398 => (x"c2",x"87",x"ed",x"c0"),
  2399 => (x"48",x"bf",x"d8",x"f5"),
  2400 => (x"03",x"a8",x"b7",x"c7"),
  2401 => (x"c2",x"87",x"c9",x"c0"),
  2402 => (x"c7",x"48",x"d8",x"f5"),
  2403 => (x"87",x"d3",x"c0",x"78"),
  2404 => (x"c1",x"48",x"66",x"c4"),
  2405 => (x"7e",x"70",x"80",x"e0"),
  2406 => (x"c0",x"02",x"bf",x"6e"),
  2407 => (x"fc",x"4b",x"87",x"c5"),
  2408 => (x"c8",x"0f",x"73",x"49"),
  2409 => (x"78",x"c1",x"48",x"a6"),
  2410 => (x"f5",x"c2",x"7e",x"c0"),
  2411 => (x"50",x"c0",x"48",x"d0"),
  2412 => (x"c3",x"49",x"ee",x"cb"),
  2413 => (x"a6",x"d4",x"87",x"c6"),
  2414 => (x"d0",x"f5",x"c2",x"58"),
  2415 => (x"c1",x"05",x"bf",x"97"),
  2416 => (x"49",x"74",x"87",x"de"),
  2417 => (x"05",x"99",x"f0",x"c3"),
  2418 => (x"c1",x"87",x"cd",x"c0"),
  2419 => (x"df",x"ff",x"49",x"da"),
  2420 => (x"98",x"70",x"87",x"c5"),
  2421 => (x"87",x"c8",x"c1",x"02"),
  2422 => (x"bf",x"e8",x"7e",x"c1"),
  2423 => (x"ff",x"c3",x"49",x"4b"),
  2424 => (x"2b",x"b7",x"c8",x"99"),
  2425 => (x"d9",x"c2",x"b3",x"71"),
  2426 => (x"ff",x"49",x"bf",x"f8"),
  2427 => (x"d0",x"87",x"e6",x"da"),
  2428 => (x"d3",x"c2",x"49",x"66"),
  2429 => (x"02",x"98",x"70",x"87"),
  2430 => (x"c2",x"87",x"c6",x"c0"),
  2431 => (x"c1",x"48",x"d0",x"f5"),
  2432 => (x"d0",x"f5",x"c2",x"50"),
  2433 => (x"c0",x"05",x"bf",x"97"),
  2434 => (x"49",x"73",x"87",x"d6"),
  2435 => (x"05",x"99",x"f0",x"c3"),
  2436 => (x"c1",x"87",x"c5",x"ff"),
  2437 => (x"dd",x"ff",x"49",x"da"),
  2438 => (x"98",x"70",x"87",x"fd"),
  2439 => (x"87",x"f8",x"fe",x"05"),
  2440 => (x"e0",x"c0",x"02",x"6e"),
  2441 => (x"48",x"a6",x"cc",x"87"),
  2442 => (x"bf",x"d8",x"f5",x"c2"),
  2443 => (x"49",x"66",x"cc",x"78"),
  2444 => (x"66",x"c4",x"91",x"cc"),
  2445 => (x"70",x"80",x"71",x"48"),
  2446 => (x"02",x"bf",x"6e",x"7e"),
  2447 => (x"4b",x"87",x"c6",x"c0"),
  2448 => (x"73",x"49",x"66",x"cc"),
  2449 => (x"02",x"66",x"c8",x"0f"),
  2450 => (x"c2",x"87",x"c8",x"c0"),
  2451 => (x"49",x"bf",x"d8",x"f5"),
  2452 => (x"ec",x"87",x"e9",x"f1"),
  2453 => (x"26",x"4d",x"26",x"8e"),
  2454 => (x"26",x"4b",x"26",x"4c"),
  2455 => (x"00",x"00",x"00",x"4f"),
  2456 => (x"00",x"00",x"00",x"00"),
  2457 => (x"14",x"11",x"12",x"58"),
  2458 => (x"23",x"1c",x"1b",x"1d"),
  2459 => (x"94",x"91",x"59",x"5a"),
  2460 => (x"f4",x"eb",x"f2",x"f5"),
  2461 => (x"00",x"00",x"00",x"00"),
  2462 => (x"00",x"00",x"00",x"00"),
  2463 => (x"ff",x"4a",x"71",x"1e"),
  2464 => (x"72",x"49",x"bf",x"c8"),
  2465 => (x"4f",x"26",x"48",x"a1"),
  2466 => (x"bf",x"c8",x"ff",x"1e"),
  2467 => (x"c0",x"c0",x"fe",x"89"),
  2468 => (x"a9",x"c0",x"c0",x"c0"),
  2469 => (x"c0",x"87",x"c4",x"01"),
  2470 => (x"c1",x"87",x"c2",x"4a"),
  2471 => (x"26",x"48",x"72",x"4a"),
  2472 => (x"5b",x"5e",x"0e",x"4f"),
  2473 => (x"71",x"0e",x"5d",x"5c"),
  2474 => (x"4c",x"d4",x"ff",x"4b"),
  2475 => (x"c0",x"48",x"66",x"d0"),
  2476 => (x"ff",x"49",x"d6",x"78"),
  2477 => (x"c3",x"87",x"dd",x"dd"),
  2478 => (x"49",x"6c",x"7c",x"ff"),
  2479 => (x"71",x"99",x"ff",x"c3"),
  2480 => (x"f0",x"c3",x"49",x"4d"),
  2481 => (x"a9",x"e0",x"c1",x"99"),
  2482 => (x"c3",x"87",x"cb",x"05"),
  2483 => (x"48",x"6c",x"7c",x"ff"),
  2484 => (x"66",x"d0",x"98",x"c3"),
  2485 => (x"ff",x"c3",x"78",x"08"),
  2486 => (x"49",x"4a",x"6c",x"7c"),
  2487 => (x"ff",x"c3",x"31",x"c8"),
  2488 => (x"71",x"4a",x"6c",x"7c"),
  2489 => (x"c8",x"49",x"72",x"b2"),
  2490 => (x"7c",x"ff",x"c3",x"31"),
  2491 => (x"b2",x"71",x"4a",x"6c"),
  2492 => (x"31",x"c8",x"49",x"72"),
  2493 => (x"6c",x"7c",x"ff",x"c3"),
  2494 => (x"ff",x"b2",x"71",x"4a"),
  2495 => (x"e0",x"c0",x"48",x"d0"),
  2496 => (x"02",x"9b",x"73",x"78"),
  2497 => (x"7b",x"72",x"87",x"c2"),
  2498 => (x"4d",x"26",x"48",x"75"),
  2499 => (x"4b",x"26",x"4c",x"26"),
  2500 => (x"26",x"1e",x"4f",x"26"),
  2501 => (x"5b",x"5e",x"0e",x"4f"),
  2502 => (x"86",x"f8",x"0e",x"5c"),
  2503 => (x"a6",x"c8",x"1e",x"76"),
  2504 => (x"87",x"fd",x"fd",x"49"),
  2505 => (x"4b",x"70",x"86",x"c4"),
  2506 => (x"a8",x"c2",x"48",x"6e"),
  2507 => (x"87",x"f0",x"c2",x"03"),
  2508 => (x"f0",x"c3",x"4a",x"73"),
  2509 => (x"aa",x"d0",x"c1",x"9a"),
  2510 => (x"c1",x"87",x"c7",x"02"),
  2511 => (x"c2",x"05",x"aa",x"e0"),
  2512 => (x"49",x"73",x"87",x"de"),
  2513 => (x"c3",x"02",x"99",x"c8"),
  2514 => (x"87",x"c6",x"ff",x"87"),
  2515 => (x"9c",x"c3",x"4c",x"73"),
  2516 => (x"c1",x"05",x"ac",x"c2"),
  2517 => (x"66",x"c4",x"87",x"c2"),
  2518 => (x"71",x"31",x"c9",x"49"),
  2519 => (x"4a",x"66",x"c4",x"1e"),
  2520 => (x"f5",x"c2",x"92",x"d4"),
  2521 => (x"81",x"72",x"49",x"dc"),
  2522 => (x"87",x"e8",x"cd",x"fe"),
  2523 => (x"da",x"ff",x"49",x"d8"),
  2524 => (x"c0",x"c8",x"87",x"e2"),
  2525 => (x"f4",x"e3",x"c2",x"1e"),
  2526 => (x"da",x"e7",x"fd",x"49"),
  2527 => (x"48",x"d0",x"ff",x"87"),
  2528 => (x"c2",x"78",x"e0",x"c0"),
  2529 => (x"cc",x"1e",x"f4",x"e3"),
  2530 => (x"92",x"d4",x"4a",x"66"),
  2531 => (x"49",x"dc",x"f5",x"c2"),
  2532 => (x"cb",x"fe",x"81",x"72"),
  2533 => (x"86",x"cc",x"87",x"ef"),
  2534 => (x"c1",x"05",x"ac",x"c1"),
  2535 => (x"66",x"c4",x"87",x"c2"),
  2536 => (x"71",x"31",x"c9",x"49"),
  2537 => (x"4a",x"66",x"c4",x"1e"),
  2538 => (x"f5",x"c2",x"92",x"d4"),
  2539 => (x"81",x"72",x"49",x"dc"),
  2540 => (x"87",x"e0",x"cc",x"fe"),
  2541 => (x"1e",x"f4",x"e3",x"c2"),
  2542 => (x"d4",x"4a",x"66",x"c8"),
  2543 => (x"dc",x"f5",x"c2",x"92"),
  2544 => (x"fe",x"81",x"72",x"49"),
  2545 => (x"d7",x"87",x"ef",x"c9"),
  2546 => (x"c7",x"d9",x"ff",x"49"),
  2547 => (x"1e",x"c0",x"c8",x"87"),
  2548 => (x"49",x"f4",x"e3",x"c2"),
  2549 => (x"87",x"dc",x"e5",x"fd"),
  2550 => (x"d0",x"ff",x"86",x"cc"),
  2551 => (x"78",x"e0",x"c0",x"48"),
  2552 => (x"4c",x"26",x"8e",x"f8"),
  2553 => (x"4f",x"26",x"4b",x"26"),
  2554 => (x"5c",x"5b",x"5e",x"0e"),
  2555 => (x"86",x"fc",x"0e",x"5d"),
  2556 => (x"d4",x"ff",x"4d",x"71"),
  2557 => (x"7e",x"66",x"d4",x"4c"),
  2558 => (x"a8",x"b7",x"c3",x"48"),
  2559 => (x"87",x"e2",x"c1",x"01"),
  2560 => (x"66",x"c4",x"1e",x"75"),
  2561 => (x"c2",x"93",x"d4",x"4b"),
  2562 => (x"73",x"83",x"dc",x"f5"),
  2563 => (x"e4",x"c3",x"fe",x"49"),
  2564 => (x"49",x"a3",x"c8",x"87"),
  2565 => (x"d0",x"ff",x"49",x"69"),
  2566 => (x"78",x"e1",x"c8",x"48"),
  2567 => (x"48",x"71",x"7c",x"dd"),
  2568 => (x"70",x"98",x"ff",x"c3"),
  2569 => (x"c8",x"4a",x"71",x"7c"),
  2570 => (x"48",x"72",x"2a",x"b7"),
  2571 => (x"70",x"98",x"ff",x"c3"),
  2572 => (x"d0",x"4a",x"71",x"7c"),
  2573 => (x"48",x"72",x"2a",x"b7"),
  2574 => (x"70",x"98",x"ff",x"c3"),
  2575 => (x"d8",x"48",x"71",x"7c"),
  2576 => (x"7c",x"70",x"28",x"b7"),
  2577 => (x"7c",x"7c",x"7c",x"c0"),
  2578 => (x"7c",x"7c",x"7c",x"7c"),
  2579 => (x"7c",x"7c",x"7c",x"7c"),
  2580 => (x"48",x"d0",x"ff",x"7c"),
  2581 => (x"c4",x"78",x"e0",x"c0"),
  2582 => (x"49",x"dc",x"1e",x"66"),
  2583 => (x"87",x"d9",x"d7",x"ff"),
  2584 => (x"8e",x"fc",x"86",x"c8"),
  2585 => (x"4c",x"26",x"4d",x"26"),
  2586 => (x"4f",x"26",x"4b",x"26"),
  2587 => (x"c0",x"1e",x"73",x"1e"),
  2588 => (x"e2",x"c2",x"1e",x"4b"),
  2589 => (x"fd",x"49",x"bf",x"e8"),
  2590 => (x"86",x"c4",x"87",x"ee"),
  2591 => (x"bf",x"ec",x"e2",x"c2"),
  2592 => (x"c1",x"dc",x"fe",x"49"),
  2593 => (x"05",x"98",x"70",x"87"),
  2594 => (x"e2",x"c2",x"87",x"c4"),
  2595 => (x"48",x"73",x"4b",x"d4"),
  2596 => (x"4f",x"26",x"4b",x"26"),
  2597 => (x"20",x"4d",x"4f",x"52"),
  2598 => (x"64",x"61",x"6f",x"6c"),
  2599 => (x"20",x"67",x"6e",x"69"),
  2600 => (x"6c",x"69",x"61",x"66"),
  2601 => (x"00",x"00",x"64",x"65"),
  2602 => (x"00",x"00",x"28",x"b0"),
  2603 => (x"00",x"00",x"28",x"bc"),
  2604 => (x"20",x"43",x"42",x"42"),
  2605 => (x"20",x"20",x"20",x"20"),
  2606 => (x"00",x"44",x"48",x"56"),
  2607 => (x"20",x"43",x"42",x"42"),
  2608 => (x"20",x"20",x"20",x"20"),
  2609 => (x"00",x"4d",x"4f",x"52"),
  2610 => (x"00",x"00",x"1b",x"ab"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

