library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"7c40407c",
     1 => x"1c00007c",
     2 => x"3c60603c",
     3 => x"7c3c001c",
     4 => x"7c603060",
     5 => x"6c44003c",
     6 => x"6c381038",
     7 => x"1c000044",
     8 => x"3c60e0bc",
     9 => x"4400001c",
    10 => x"4c5c7464",
    11 => x"08000044",
    12 => x"41773e08",
    13 => x"00000041",
    14 => x"007f7f00",
    15 => x"41000000",
    16 => x"083e7741",
    17 => x"01020008",
    18 => x"02020301",
    19 => x"7f7f0001",
    20 => x"7f7f7f7f",
    21 => x"0808007f",
    22 => x"3e3e1c1c",
    23 => x"7f7f7f7f",
    24 => x"1c1c3e3e",
    25 => x"10000808",
    26 => x"187c7c18",
    27 => x"10000010",
    28 => x"307c7c30",
    29 => x"30100010",
    30 => x"1e786060",
    31 => x"66420006",
    32 => x"663c183c",
    33 => x"38780042",
    34 => x"6cc6c26a",
    35 => x"00600038",
    36 => x"00006000",
    37 => x"5e0e0060",
    38 => x"0e5d5c5b",
    39 => x"c24c711e",
    40 => x"4dbfd9ee",
    41 => x"1ec04bc0",
    42 => x"c702ab74",
    43 => x"48a6c487",
    44 => x"87c578c0",
    45 => x"c148a6c4",
    46 => x"1e66c478",
    47 => x"dfee4973",
    48 => x"c086c887",
    49 => x"eeef49e0",
    50 => x"4aa5c487",
    51 => x"f0f0496a",
    52 => x"87c6f187",
    53 => x"83c185cb",
    54 => x"04abb7c8",
    55 => x"2687c7ff",
    56 => x"4c264d26",
    57 => x"4f264b26",
    58 => x"c24a711e",
    59 => x"c25addee",
    60 => x"c748ddee",
    61 => x"ddfe4978",
    62 => x"1e4f2687",
    63 => x"4a711e73",
    64 => x"03aab7c0",
    65 => x"d2c287d3",
    66 => x"c405bffe",
    67 => x"c24bc187",
    68 => x"c24bc087",
    69 => x"c45bc2d3",
    70 => x"c2d3c287",
    71 => x"fed2c25a",
    72 => x"9ac14abf",
    73 => x"49a2c0c1",
    74 => x"fc87e8ec",
    75 => x"fed2c248",
    76 => x"effe78bf",
    77 => x"4a711e87",
    78 => x"721e66c4",
    79 => x"87f9ea49",
    80 => x"1e4f2626",
    81 => x"c348d4ff",
    82 => x"d0ff78ff",
    83 => x"78e1c048",
    84 => x"c148d4ff",
    85 => x"c4487178",
    86 => x"08d4ff30",
    87 => x"48d0ff78",
    88 => x"2678e0c0",
    89 => x"d2c21e4f",
    90 => x"e649bffe",
    91 => x"eec287f9",
    92 => x"bfe848d1",
    93 => x"cdeec278",
    94 => x"78bfec48",
    95 => x"bfd1eec2",
    96 => x"ffc3494a",
    97 => x"2ab7c899",
    98 => x"b0714872",
    99 => x"58d9eec2",
   100 => x"5e0e4f26",
   101 => x"0e5d5c5b",
   102 => x"c8ff4b71",
   103 => x"cceec287",
   104 => x"7350c048",
   105 => x"87dfe649",
   106 => x"c24c4970",
   107 => x"49eecb9c",
   108 => x"7087d3cc",
   109 => x"cceec24d",
   110 => x"c105bf97",
   111 => x"66d087e2",
   112 => x"d5eec249",
   113 => x"d60599bf",
   114 => x"4966d487",
   115 => x"bfcdeec2",
   116 => x"87cb0599",
   117 => x"eee54973",
   118 => x"02987087",
   119 => x"c187c1c1",
   120 => x"87c1fe4c",
   121 => x"e9cb4975",
   122 => x"02987087",
   123 => x"eec287c6",
   124 => x"50c148cc",
   125 => x"97cceec2",
   126 => x"e3c005bf",
   127 => x"d5eec287",
   128 => x"66d049bf",
   129 => x"d6ff0599",
   130 => x"cdeec287",
   131 => x"66d449bf",
   132 => x"caff0599",
   133 => x"e4497387",
   134 => x"987087ed",
   135 => x"87fffe05",
   136 => x"fbfa4874",
   137 => x"5b5e0e87",
   138 => x"f80e5d5c",
   139 => x"4c4dc086",
   140 => x"c47ebfec",
   141 => x"eec248a6",
   142 => x"c178bfd9",
   143 => x"c71ec01e",
   144 => x"87cefd49",
   145 => x"987086c8",
   146 => x"ff87cd02",
   147 => x"87ebfa49",
   148 => x"e349dac1",
   149 => x"4dc187f1",
   150 => x"97cceec2",
   151 => x"87cf02bf",
   152 => x"bfe6d2c2",
   153 => x"c2b9c149",
   154 => x"7159ead2",
   155 => x"c287d4fb",
   156 => x"4bbfd1ee",
   157 => x"bffed2c2",
   158 => x"87d9c105",
   159 => x"c848a6c4",
   160 => x"c278c0c0",
   161 => x"6e7eead2",
   162 => x"6e49bf97",
   163 => x"7080c148",
   164 => x"f2e2717e",
   165 => x"02987087",
   166 => x"66c487c3",
   167 => x"4866c4b3",
   168 => x"c828b7c1",
   169 => x"987058a6",
   170 => x"87dbff05",
   171 => x"e249fdc3",
   172 => x"fac387d5",
   173 => x"87cfe249",
   174 => x"ffc34973",
   175 => x"c01e7199",
   176 => x"87f1f949",
   177 => x"b7c84973",
   178 => x"c11e7129",
   179 => x"87e5f949",
   180 => x"fac586c8",
   181 => x"d5eec287",
   182 => x"029b4bbf",
   183 => x"d2c287dd",
   184 => x"c749bffa",
   185 => x"987087ec",
   186 => x"c087c405",
   187 => x"c287d24b",
   188 => x"d1c749e0",
   189 => x"fed2c287",
   190 => x"c287c658",
   191 => x"c048fad2",
   192 => x"c2497378",
   193 => x"87ce0599",
   194 => x"e049ebc3",
   195 => x"497087f9",
   196 => x"c00299c2",
   197 => x"4cfb87c2",
   198 => x"99c14973",
   199 => x"c387ce05",
   200 => x"e2e049f4",
   201 => x"c2497087",
   202 => x"c2c00299",
   203 => x"734cfa87",
   204 => x"0599c849",
   205 => x"f5c387cd",
   206 => x"87cbe049",
   207 => x"99c24970",
   208 => x"c287d602",
   209 => x"02bfddee",
   210 => x"4887cac0",
   211 => x"eec288c1",
   212 => x"c2c058e1",
   213 => x"c14cff87",
   214 => x"c449734d",
   215 => x"cec00599",
   216 => x"49f2c387",
   217 => x"87dfdfff",
   218 => x"99c24970",
   219 => x"c287dc02",
   220 => x"7ebfddee",
   221 => x"a8b7c748",
   222 => x"87cbc003",
   223 => x"80c1486e",
   224 => x"58e1eec2",
   225 => x"fe87c2c0",
   226 => x"c34dc14c",
   227 => x"deff49fd",
   228 => x"497087f5",
   229 => x"c00299c2",
   230 => x"eec287d5",
   231 => x"c002bfdd",
   232 => x"eec287c9",
   233 => x"78c048dd",
   234 => x"fd87c2c0",
   235 => x"c34dc14c",
   236 => x"deff49fa",
   237 => x"497087d1",
   238 => x"c00299c2",
   239 => x"eec287d9",
   240 => x"c748bfdd",
   241 => x"c003a8b7",
   242 => x"eec287c9",
   243 => x"78c748dd",
   244 => x"fc87c2c0",
   245 => x"c04dc14c",
   246 => x"c003acb7",
   247 => x"66c487d3",
   248 => x"80d8c148",
   249 => x"bf6e7e70",
   250 => x"87c5c002",
   251 => x"7349744b",
   252 => x"c31ec00f",
   253 => x"dac11ef0",
   254 => x"87d6f649",
   255 => x"987086c8",
   256 => x"87d8c002",
   257 => x"bfddeec2",
   258 => x"cb496e7e",
   259 => x"4a66c491",
   260 => x"026a8271",
   261 => x"4b87c5c0",
   262 => x"0f73496e",
   263 => x"c0029d75",
   264 => x"eec287c8",
   265 => x"f149bfdd",
   266 => x"d3c287ec",
   267 => x"c002bfc2",
   268 => x"c24987dd",
   269 => x"987087dc",
   270 => x"87d3c002",
   271 => x"bfddeec2",
   272 => x"87d2f149",
   273 => x"f2f249c0",
   274 => x"c2d3c287",
   275 => x"f878c048",
   276 => x"87ccf28e",
   277 => x"5c5b5e0e",
   278 => x"711e0e5d",
   279 => x"d9eec24c",
   280 => x"cdc149bf",
   281 => x"d1c14da1",
   282 => x"747e6981",
   283 => x"87cf029c",
   284 => x"744ba5c4",
   285 => x"d9eec27b",
   286 => x"ebf149bf",
   287 => x"747b6e87",
   288 => x"87c4059c",
   289 => x"87c24bc0",
   290 => x"49734bc1",
   291 => x"d487ecf1",
   292 => x"87c80266",
   293 => x"87eec049",
   294 => x"87c24a70",
   295 => x"d3c24ac0",
   296 => x"f0265ac6",
   297 => x"000087fa",
   298 => x"12580000",
   299 => x"1b1d1411",
   300 => x"595a231c",
   301 => x"f2f59491",
   302 => x"0000f4eb",
   303 => x"00000000",
   304 => x"00000000",
   305 => x"711e0000",
   306 => x"bfc8ff4a",
   307 => x"48a17249",
   308 => x"ff1e4f26",
   309 => x"fe89bfc8",
   310 => x"c0c0c0c0",
   311 => x"c401a9c0",
   312 => x"c24ac087",
   313 => x"724ac187",
   314 => x"0e4f2648",
   315 => x"5d5c5b5e",
   316 => x"ff4b710e",
   317 => x"66d04cd4",
   318 => x"d678c048",
   319 => x"fedaff49",
   320 => x"7cffc387",
   321 => x"ffc3496c",
   322 => x"494d7199",
   323 => x"c199f0c3",
   324 => x"cb05a9e0",
   325 => x"7cffc387",
   326 => x"98c3486c",
   327 => x"780866d0",
   328 => x"6c7cffc3",
   329 => x"31c8494a",
   330 => x"6c7cffc3",
   331 => x"72b2714a",
   332 => x"c331c849",
   333 => x"4a6c7cff",
   334 => x"4972b271",
   335 => x"ffc331c8",
   336 => x"714a6c7c",
   337 => x"48d0ffb2",
   338 => x"7378e0c0",
   339 => x"87c2029b",
   340 => x"48757b72",
   341 => x"4c264d26",
   342 => x"4f264b26",
   343 => x"0e4f261e",
   344 => x"0e5c5b5e",
   345 => x"1e7686f8",
   346 => x"fd49a6c8",
   347 => x"86c487fd",
   348 => x"486e4b70",
   349 => x"c203a8c2",
   350 => x"4a7387f0",
   351 => x"c19af0c3",
   352 => x"c702aad0",
   353 => x"aae0c187",
   354 => x"87dec205",
   355 => x"99c84973",
   356 => x"ff87c302",
   357 => x"4c7387c6",
   358 => x"acc29cc3",
   359 => x"87c2c105",
   360 => x"c94966c4",
   361 => x"c41e7131",
   362 => x"92d44a66",
   363 => x"49e1eec2",
   364 => x"d0fe8172",
   365 => x"49d887d1",
   366 => x"87c3d8ff",
   367 => x"c21ec0c8",
   368 => x"fd49fedc",
   369 => x"ff87d7ec",
   370 => x"e0c048d0",
   371 => x"fedcc278",
   372 => x"4a66cc1e",
   373 => x"eec292d4",
   374 => x"817249e1",
   375 => x"87d9cefe",
   376 => x"acc186cc",
   377 => x"87c2c105",
   378 => x"c94966c4",
   379 => x"c41e7131",
   380 => x"92d44a66",
   381 => x"49e1eec2",
   382 => x"cffe8172",
   383 => x"dcc287c9",
   384 => x"66c81efe",
   385 => x"c292d44a",
   386 => x"7249e1ee",
   387 => x"daccfe81",
   388 => x"ff49d787",
   389 => x"c887e8d6",
   390 => x"dcc21ec0",
   391 => x"eafd49fe",
   392 => x"86cc87d5",
   393 => x"c048d0ff",
   394 => x"8ef878e0",
   395 => x"0e87e7fc",
   396 => x"5d5c5b5e",
   397 => x"4d711e0e",
   398 => x"d44cd4ff",
   399 => x"c3487e66",
   400 => x"c506a8b7",
   401 => x"c148c087",
   402 => x"497587e9",
   403 => x"87ffdcfe",
   404 => x"66c41e75",
   405 => x"c293d44b",
   406 => x"7383e1ee",
   407 => x"d8c6fe49",
   408 => x"6b83c887",
   409 => x"48d0ff4b",
   410 => x"dd78e1c8",
   411 => x"c348737c",
   412 => x"7c7098ff",
   413 => x"b7c84973",
   414 => x"c3487129",
   415 => x"7c7098ff",
   416 => x"b7d04973",
   417 => x"c3487129",
   418 => x"7c7098ff",
   419 => x"b7d84873",
   420 => x"c07c7028",
   421 => x"7c7c7c7c",
   422 => x"7c7c7c7c",
   423 => x"7c7c7c7c",
   424 => x"c048d0ff",
   425 => x"66c478e0",
   426 => x"ff49dc1e",
   427 => x"c887f5d4",
   428 => x"26487386",
   429 => x"1e87ddfa",
   430 => x"4bc01e73",
   431 => x"f8dbc21e",
   432 => x"eafd49bf",
   433 => x"c286c487",
   434 => x"49bffcdb",
   435 => x"87e3defe",
   436 => x"c4059870",
   437 => x"e5dbc287",
   438 => x"c448734b",
   439 => x"264d2687",
   440 => x"264b264c",
   441 => x"4d4f524f",
   442 => x"616f6c20",
   443 => x"676e6964",
   444 => x"69616620",
   445 => x"0064656c",
   446 => x"00002700",
   447 => x"0000270c",
   448 => x"20434242",
   449 => x"20202020",
   450 => x"00444856",
   451 => x"20434242",
   452 => x"20202020",
   453 => x"004d4f52",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
