library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f0f4c287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49f0f4c2",
    18 => x"48f8e1c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"f8e1c287",
    25 => x"f4e1c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e8c187f7",
    29 => x"e1c287c6",
    30 => x"e1c24df8",
    31 => x"ad744cf8",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"731e741e",
    65 => x"c11e721e",
    66 => x"87d0048b",
    67 => x"02114812",
    68 => x"c34c87ca",
    69 => x"749c98df",
    70 => x"87eb0288",
    71 => x"4b264a26",
    72 => x"4f264c26",
    73 => x"8148731e",
    74 => x"c502a973",
    75 => x"05531287",
    76 => x"4f2687f6",
    77 => x"711e731e",
    78 => x"4b66c84a",
    79 => x"718bc149",
    80 => x"87cf0299",
    81 => x"d4ff4812",
    82 => x"49737808",
    83 => x"99718bc1",
    84 => x"2687f105",
    85 => x"0e4f264b",
    86 => x"0e5c5b5e",
    87 => x"d4ff4a71",
    88 => x"4b66cc4c",
    89 => x"718bc149",
    90 => x"87ce0299",
    91 => x"6c7cffc3",
    92 => x"c1497352",
    93 => x"0599718b",
    94 => x"4c2687f2",
    95 => x"4f264b26",
    96 => x"ff1e731e",
    97 => x"ffc34bd4",
    98 => x"c34a6b7b",
    99 => x"496b7bff",
   100 => x"b17232c8",
   101 => x"6b7bffc3",
   102 => x"7131c84a",
   103 => x"7bffc3b2",
   104 => x"32c8496b",
   105 => x"4871b172",
   106 => x"4f264b26",
   107 => x"5c5b5e0e",
   108 => x"4d710e5d",
   109 => x"754cd4ff",
   110 => x"98ffc348",
   111 => x"e1c27c70",
   112 => x"c805bff8",
   113 => x"4866d087",
   114 => x"a6d430c9",
   115 => x"4966d058",
   116 => x"487129d8",
   117 => x"7098ffc3",
   118 => x"4966d07c",
   119 => x"487129d0",
   120 => x"7098ffc3",
   121 => x"4966d07c",
   122 => x"487129c8",
   123 => x"7098ffc3",
   124 => x"4866d07c",
   125 => x"7098ffc3",
   126 => x"d049757c",
   127 => x"c3487129",
   128 => x"7c7098ff",
   129 => x"f0c94b6c",
   130 => x"ffc34aff",
   131 => x"87cf05ab",
   132 => x"6c7c7149",
   133 => x"028ac14b",
   134 => x"ab7187c5",
   135 => x"7387f202",
   136 => x"264d2648",
   137 => x"264b264c",
   138 => x"49c01e4f",
   139 => x"c348d4ff",
   140 => x"81c178ff",
   141 => x"a9b7c8c3",
   142 => x"2687f104",
   143 => x"5b5e0e4f",
   144 => x"c00e5d5c",
   145 => x"f7c1f0ff",
   146 => x"c0c0c14d",
   147 => x"4bc0c0c0",
   148 => x"c487d6ff",
   149 => x"c04cdff8",
   150 => x"fd49751e",
   151 => x"86c487ce",
   152 => x"c005a8c1",
   153 => x"d4ff87e5",
   154 => x"78ffc348",
   155 => x"e1c01e73",
   156 => x"49e9c1f0",
   157 => x"c487f5fc",
   158 => x"05987086",
   159 => x"d4ff87ca",
   160 => x"78ffc348",
   161 => x"87cb48c1",
   162 => x"c187defe",
   163 => x"c6ff058c",
   164 => x"2648c087",
   165 => x"264c264d",
   166 => x"0e4f264b",
   167 => x"0e5c5b5e",
   168 => x"c1f0ffc0",
   169 => x"d4ff4cc1",
   170 => x"78ffc348",
   171 => x"f749e0cb",
   172 => x"4bd387f5",
   173 => x"49741ec0",
   174 => x"c487f1fb",
   175 => x"05987086",
   176 => x"d4ff87ca",
   177 => x"78ffc348",
   178 => x"87cb48c1",
   179 => x"c187dafd",
   180 => x"dfff058b",
   181 => x"2648c087",
   182 => x"264b264c",
   183 => x"0000004f",
   184 => x"00444d43",
   185 => x"5c5b5e0e",
   186 => x"ffc30e5d",
   187 => x"4bd4ff4d",
   188 => x"c687f6fc",
   189 => x"e1c01eea",
   190 => x"49c8c1f0",
   191 => x"c487edfa",
   192 => x"02a8c186",
   193 => x"d2fe87c8",
   194 => x"c148c087",
   195 => x"eff987e8",
   196 => x"cf497087",
   197 => x"c699ffff",
   198 => x"c802a9ea",
   199 => x"87fbfd87",
   200 => x"d1c148c0",
   201 => x"c07b7587",
   202 => x"d0fc4cf1",
   203 => x"02987087",
   204 => x"c087ecc0",
   205 => x"f0ffc01e",
   206 => x"f949fac1",
   207 => x"86c487ee",
   208 => x"da059870",
   209 => x"6b7b7587",
   210 => x"757b7549",
   211 => x"757b757b",
   212 => x"99c0c17b",
   213 => x"c187c402",
   214 => x"c087db48",
   215 => x"c287d748",
   216 => x"87ca05ac",
   217 => x"f449c0ce",
   218 => x"48c087fd",
   219 => x"8cc187c8",
   220 => x"87f6fe05",
   221 => x"4d2648c0",
   222 => x"4b264c26",
   223 => x"00004f26",
   224 => x"43484453",
   225 => x"69616620",
   226 => x"000a216c",
   227 => x"5c5b5e0e",
   228 => x"d0ff0e5d",
   229 => x"d0e5c04d",
   230 => x"c24cc0c1",
   231 => x"c148f8e1",
   232 => x"49d8d078",
   233 => x"c787c0f4",
   234 => x"f97dc24b",
   235 => x"7dc387fb",
   236 => x"49741ec0",
   237 => x"c487f5f7",
   238 => x"05a8c186",
   239 => x"c24b87c1",
   240 => x"87cb05ab",
   241 => x"f349d0d0",
   242 => x"48c087dd",
   243 => x"c187f6c0",
   244 => x"d4ff058b",
   245 => x"87ccfc87",
   246 => x"58fce1c2",
   247 => x"cd059870",
   248 => x"c01ec187",
   249 => x"d0c1f0ff",
   250 => x"87c0f749",
   251 => x"d4ff86c4",
   252 => x"78ffc348",
   253 => x"c287ccc5",
   254 => x"c258c0e2",
   255 => x"48d4ff7d",
   256 => x"c178ffc3",
   257 => x"264d2648",
   258 => x"264b264c",
   259 => x"0000004f",
   260 => x"52524549",
   261 => x"00000000",
   262 => x"00495053",
   263 => x"5c5b5e0e",
   264 => x"4d710e5d",
   265 => x"ff4cffc3",
   266 => x"7b744bd4",
   267 => x"c448d0ff",
   268 => x"7b7478c3",
   269 => x"ffc01e75",
   270 => x"49d8c1f0",
   271 => x"c487edf5",
   272 => x"02987086",
   273 => x"c8d287cb",
   274 => x"87dbf149",
   275 => x"eec048c1",
   276 => x"c37b7487",
   277 => x"c0c87bfe",
   278 => x"4966d41e",
   279 => x"c487d5f3",
   280 => x"747b7486",
   281 => x"d87b747b",
   282 => x"744ae0da",
   283 => x"c5056b7b",
   284 => x"058ac187",
   285 => x"7b7487f5",
   286 => x"c248d0ff",
   287 => x"2648c078",
   288 => x"264c264d",
   289 => x"004f264b",
   290 => x"74697257",
   291 => x"61662065",
   292 => x"64656c69",
   293 => x"5e0e000a",
   294 => x"0e5d5c5b",
   295 => x"4b7186fc",
   296 => x"c04cd4ff",
   297 => x"cdeec57e",
   298 => x"ffc34adf",
   299 => x"c3486c7c",
   300 => x"c005a8fe",
   301 => x"4d7487f8",
   302 => x"cc029b73",
   303 => x"1e66d487",
   304 => x"d2f24973",
   305 => x"d486c487",
   306 => x"48d0ff87",
   307 => x"d478d1c4",
   308 => x"ffc34a66",
   309 => x"058ac17d",
   310 => x"a6d887f8",
   311 => x"7cffc35a",
   312 => x"059b737c",
   313 => x"d0ff87c5",
   314 => x"c178d048",
   315 => x"8ac17e4a",
   316 => x"87f6fe05",
   317 => x"8efc486e",
   318 => x"4c264d26",
   319 => x"4f264b26",
   320 => x"711e731e",
   321 => x"ff4bc04a",
   322 => x"ffc348d4",
   323 => x"48d0ff78",
   324 => x"ff78c3c4",
   325 => x"ffc348d4",
   326 => x"c01e7278",
   327 => x"d1c1f0ff",
   328 => x"87c8f249",
   329 => x"987086c4",
   330 => x"c887d205",
   331 => x"66cc1ec0",
   332 => x"87e2fd49",
   333 => x"4b7086c4",
   334 => x"c248d0ff",
   335 => x"26487378",
   336 => x"0e4f264b",
   337 => x"5d5c5b5e",
   338 => x"c01ec00e",
   339 => x"c9c1f0ff",
   340 => x"87d8f149",
   341 => x"e2c21ed2",
   342 => x"f9fc49c0",
   343 => x"c086c887",
   344 => x"d284c14c",
   345 => x"f804acb7",
   346 => x"c0e2c287",
   347 => x"c349bf97",
   348 => x"c0c199c0",
   349 => x"e7c005a9",
   350 => x"c7e2c287",
   351 => x"d049bf97",
   352 => x"c8e2c231",
   353 => x"c84abf97",
   354 => x"c2b17232",
   355 => x"bf97c9e2",
   356 => x"4c71b14a",
   357 => x"ffffffcf",
   358 => x"ca84c19c",
   359 => x"87e7c134",
   360 => x"97c9e2c2",
   361 => x"31c149bf",
   362 => x"e2c299c6",
   363 => x"4abf97ca",
   364 => x"722ab7c7",
   365 => x"c5e2c2b1",
   366 => x"4d4abf97",
   367 => x"e2c29dcf",
   368 => x"4abf97c6",
   369 => x"32ca9ac3",
   370 => x"97c7e2c2",
   371 => x"33c24bbf",
   372 => x"e2c2b273",
   373 => x"4bbf97c8",
   374 => x"c69bc0c3",
   375 => x"b2732bb7",
   376 => x"48c181c2",
   377 => x"49703071",
   378 => x"307548c1",
   379 => x"4c724d70",
   380 => x"947184c1",
   381 => x"adb7c0c8",
   382 => x"c187cc06",
   383 => x"c82db734",
   384 => x"01adb7c0",
   385 => x"7487f4ff",
   386 => x"264d2648",
   387 => x"264b264c",
   388 => x"5b5e0e4f",
   389 => x"f80e5d5c",
   390 => x"e8eac286",
   391 => x"c278c048",
   392 => x"c01ee0e2",
   393 => x"87d8fb49",
   394 => x"987086c4",
   395 => x"c087c505",
   396 => x"87c0c948",
   397 => x"7ec14dc0",
   398 => x"bfd8f7c0",
   399 => x"d6e3c249",
   400 => x"4bc8714a",
   401 => x"7087dfea",
   402 => x"87c20598",
   403 => x"f7c07ec0",
   404 => x"c249bfd4",
   405 => x"714af2e3",
   406 => x"c9ea4bc8",
   407 => x"05987087",
   408 => x"7ec087c2",
   409 => x"fdc0026e",
   410 => x"e6e9c287",
   411 => x"eac24dbf",
   412 => x"7ebf9fde",
   413 => x"ead6c548",
   414 => x"87c705a8",
   415 => x"bfe6e9c2",
   416 => x"6e87ce4d",
   417 => x"d5e9ca48",
   418 => x"87c502a8",
   419 => x"e3c748c0",
   420 => x"e0e2c287",
   421 => x"f949751e",
   422 => x"86c487e6",
   423 => x"c5059870",
   424 => x"c748c087",
   425 => x"f7c087ce",
   426 => x"c249bfd4",
   427 => x"714af2e3",
   428 => x"f1e84bc8",
   429 => x"05987087",
   430 => x"eac287c8",
   431 => x"78c148e8",
   432 => x"f7c087da",
   433 => x"c249bfd8",
   434 => x"714ad6e3",
   435 => x"d5e84bc8",
   436 => x"02987087",
   437 => x"c087c5c0",
   438 => x"87d8c648",
   439 => x"97deeac2",
   440 => x"d5c149bf",
   441 => x"cdc005a9",
   442 => x"dfeac287",
   443 => x"c249bf97",
   444 => x"c002a9ea",
   445 => x"48c087c5",
   446 => x"c287f9c5",
   447 => x"bf97e0e2",
   448 => x"e9c3487e",
   449 => x"cec002a8",
   450 => x"c3486e87",
   451 => x"c002a8eb",
   452 => x"48c087c5",
   453 => x"c287ddc5",
   454 => x"bf97ebe2",
   455 => x"c0059949",
   456 => x"e2c287cc",
   457 => x"49bf97ec",
   458 => x"c002a9c2",
   459 => x"48c087c5",
   460 => x"c287c1c5",
   461 => x"bf97ede2",
   462 => x"e4eac248",
   463 => x"484c7058",
   464 => x"eac288c1",
   465 => x"e2c258e8",
   466 => x"49bf97ee",
   467 => x"e2c28175",
   468 => x"4abf97ef",
   469 => x"a17232c8",
   470 => x"f8eec27e",
   471 => x"c2786e48",
   472 => x"bf97f0e2",
   473 => x"58a6c848",
   474 => x"bfe8eac2",
   475 => x"87cfc202",
   476 => x"bfd4f7c0",
   477 => x"f2e3c249",
   478 => x"4bc8714a",
   479 => x"7087e7e5",
   480 => x"c5c00298",
   481 => x"c348c087",
   482 => x"eac287ea",
   483 => x"c24cbfe0",
   484 => x"c25cccef",
   485 => x"bf97c5e3",
   486 => x"c231c849",
   487 => x"bf97c4e3",
   488 => x"c249a14a",
   489 => x"bf97c6e3",
   490 => x"7232d04a",
   491 => x"e3c249a1",
   492 => x"4abf97c7",
   493 => x"a17232d8",
   494 => x"9166c449",
   495 => x"bff8eec2",
   496 => x"c0efc281",
   497 => x"cde3c259",
   498 => x"c84abf97",
   499 => x"cce3c232",
   500 => x"a24bbf97",
   501 => x"cee3c24a",
   502 => x"d04bbf97",
   503 => x"4aa27333",
   504 => x"97cfe3c2",
   505 => x"9bcf4bbf",
   506 => x"a27333d8",
   507 => x"c4efc24a",
   508 => x"748ac25a",
   509 => x"c4efc292",
   510 => x"78a17248",
   511 => x"c287c1c1",
   512 => x"bf97f2e2",
   513 => x"c231c849",
   514 => x"bf97f1e2",
   515 => x"c549a14a",
   516 => x"81ffc731",
   517 => x"efc229c9",
   518 => x"e2c259cc",
   519 => x"4abf97f7",
   520 => x"e2c232c8",
   521 => x"4bbf97f6",
   522 => x"66c44aa2",
   523 => x"c2826e92",
   524 => x"c25ac8ef",
   525 => x"c048c0ef",
   526 => x"fceec278",
   527 => x"78a17248",
   528 => x"48ccefc2",
   529 => x"bfc0efc2",
   530 => x"d0efc278",
   531 => x"c4efc248",
   532 => x"eac278bf",
   533 => x"c002bfe8",
   534 => x"487487c9",
   535 => x"7e7030c4",
   536 => x"c287c9c0",
   537 => x"48bfc8ef",
   538 => x"7e7030c4",
   539 => x"48eceac2",
   540 => x"48c1786e",
   541 => x"4d268ef8",
   542 => x"4b264c26",
   543 => x"5e0e4f26",
   544 => x"0e5d5c5b",
   545 => x"eac24a71",
   546 => x"cb02bfe8",
   547 => x"c74b7287",
   548 => x"c14d722b",
   549 => x"87c99dff",
   550 => x"2bc84b72",
   551 => x"ffc34d72",
   552 => x"f8eec29d",
   553 => x"f7c083bf",
   554 => x"02abbfd0",
   555 => x"f7c087d9",
   556 => x"e2c25bd4",
   557 => x"49731ee0",
   558 => x"c487c5f1",
   559 => x"05987086",
   560 => x"48c087c5",
   561 => x"c287e6c0",
   562 => x"02bfe8ea",
   563 => x"497587d2",
   564 => x"e2c291c4",
   565 => x"4c6981e0",
   566 => x"ffffffcf",
   567 => x"87cb9cff",
   568 => x"91c24975",
   569 => x"81e0e2c2",
   570 => x"744c699f",
   571 => x"264d2648",
   572 => x"264b264c",
   573 => x"5b5e0e4f",
   574 => x"f40e5d5c",
   575 => x"59a6cc86",
   576 => x"c50566c8",
   577 => x"c348c087",
   578 => x"66c887c7",
   579 => x"7080c848",
   580 => x"78c0487e",
   581 => x"c70266dc",
   582 => x"9766dc87",
   583 => x"87c505bf",
   584 => x"ecc248c0",
   585 => x"c11ec087",
   586 => x"e9ca4949",
   587 => x"7086c487",
   588 => x"c0029c4c",
   589 => x"eac287fc",
   590 => x"66dc4af0",
   591 => x"cadeff49",
   592 => x"02987087",
   593 => x"7487ebc0",
   594 => x"4966dc4a",
   595 => x"deff4bcb",
   596 => x"987087ee",
   597 => x"c087db02",
   598 => x"029c741e",
   599 => x"4dc087c4",
   600 => x"4dc187c2",
   601 => x"edc94975",
   602 => x"7086c487",
   603 => x"ff059c4c",
   604 => x"9c7487c4",
   605 => x"87d7c102",
   606 => x"6e49a4dc",
   607 => x"da786948",
   608 => x"66c849a4",
   609 => x"c880c448",
   610 => x"699f58a6",
   611 => x"0866c448",
   612 => x"e8eac278",
   613 => x"87d202bf",
   614 => x"9f49a4d4",
   615 => x"ffc04969",
   616 => x"487199ff",
   617 => x"7e7030d0",
   618 => x"7ec087c2",
   619 => x"66c4486e",
   620 => x"66c480bf",
   621 => x"66c87808",
   622 => x"c878c048",
   623 => x"81cc4966",
   624 => x"79bf66c4",
   625 => x"d04966c8",
   626 => x"c179c081",
   627 => x"c087c248",
   628 => x"268ef448",
   629 => x"264c264d",
   630 => x"0e4f264b",
   631 => x"5d5c5b5e",
   632 => x"d04c710e",
   633 => x"9c744d66",
   634 => x"87c2c102",
   635 => x"6949a4c8",
   636 => x"87fac002",
   637 => x"7585496c",
   638 => x"e4eac2b9",
   639 => x"baff4abf",
   640 => x"99719972",
   641 => x"87e4c002",
   642 => x"6b4ba4c4",
   643 => x"87eef949",
   644 => x"eac27b70",
   645 => x"6c49bfe0",
   646 => x"757c7181",
   647 => x"e4eac2b9",
   648 => x"baff4abf",
   649 => x"99719972",
   650 => x"87dcff05",
   651 => x"4d267c75",
   652 => x"4b264c26",
   653 => x"731e4f26",
   654 => x"9b4b711e",
   655 => x"c887c702",
   656 => x"056949a3",
   657 => x"48c087c5",
   658 => x"c287f6c0",
   659 => x"49bffcee",
   660 => x"6a4aa3c4",
   661 => x"c28ac24a",
   662 => x"92bfe0ea",
   663 => x"c249a172",
   664 => x"4abfe4ea",
   665 => x"a1729a6b",
   666 => x"d4f7c049",
   667 => x"1e66c859",
   668 => x"87ccea71",
   669 => x"987086c4",
   670 => x"c087c405",
   671 => x"c187c248",
   672 => x"264b2648",
   673 => x"1e731e4f",
   674 => x"029b4b71",
   675 => x"a3c887c7",
   676 => x"c5056949",
   677 => x"c048c087",
   678 => x"eec287f6",
   679 => x"c449bffc",
   680 => x"4a6a4aa3",
   681 => x"eac28ac2",
   682 => x"7292bfe0",
   683 => x"eac249a1",
   684 => x"6b4abfe4",
   685 => x"49a1729a",
   686 => x"59d4f7c0",
   687 => x"711e66c8",
   688 => x"c487d9e5",
   689 => x"05987086",
   690 => x"48c087c4",
   691 => x"48c187c2",
   692 => x"4f264b26",
   693 => x"5c5b5e0e",
   694 => x"86fc0e5d",
   695 => x"66d44b71",
   696 => x"029b734d",
   697 => x"c887ccc1",
   698 => x"026949a3",
   699 => x"d087c4c1",
   700 => x"eac24ca3",
   701 => x"ff49bfe4",
   702 => x"994a6cb9",
   703 => x"a966d47e",
   704 => x"c087cd06",
   705 => x"a3cc7c7b",
   706 => x"49a3c44a",
   707 => x"87ca796a",
   708 => x"c0f84972",
   709 => x"4d66d499",
   710 => x"49758d71",
   711 => x"1e7129c9",
   712 => x"f6fa4973",
   713 => x"e0e2c287",
   714 => x"fc49731e",
   715 => x"86c887c8",
   716 => x"fc7c66d4",
   717 => x"264d268e",
   718 => x"264b264c",
   719 => x"1e731e4f",
   720 => x"029b4b71",
   721 => x"c287e4c0",
   722 => x"735bd0ef",
   723 => x"c28ac24a",
   724 => x"49bfe0ea",
   725 => x"fceec292",
   726 => x"807248bf",
   727 => x"58d4efc2",
   728 => x"30c44871",
   729 => x"58f0eac2",
   730 => x"c287edc0",
   731 => x"c248ccef",
   732 => x"78bfc0ef",
   733 => x"48d0efc2",
   734 => x"bfc4efc2",
   735 => x"e8eac278",
   736 => x"87c902bf",
   737 => x"bfe0eac2",
   738 => x"c731c449",
   739 => x"c8efc287",
   740 => x"31c449bf",
   741 => x"59f0eac2",
   742 => x"4f264b26",
   743 => x"5c5b5e0e",
   744 => x"c04a710e",
   745 => x"029a724b",
   746 => x"da87e0c0",
   747 => x"699f49a2",
   748 => x"e8eac24b",
   749 => x"87cf02bf",
   750 => x"9f49a2d4",
   751 => x"c04c4969",
   752 => x"d09cffff",
   753 => x"c087c234",
   754 => x"73b3744c",
   755 => x"87edfd49",
   756 => x"4b264c26",
   757 => x"5e0e4f26",
   758 => x"0e5d5c5b",
   759 => x"a6c886f0",
   760 => x"ffffcf59",
   761 => x"c04cf8ff",
   762 => x"0266c47e",
   763 => x"e2c287d8",
   764 => x"78c048dc",
   765 => x"48d4e2c2",
   766 => x"bfd0efc2",
   767 => x"d8e2c278",
   768 => x"ccefc248",
   769 => x"eac278bf",
   770 => x"50c048fd",
   771 => x"bfeceac2",
   772 => x"dce2c249",
   773 => x"aa714abf",
   774 => x"87cbc403",
   775 => x"99cf4972",
   776 => x"87e9c005",
   777 => x"48d0f7c0",
   778 => x"bfd4e2c2",
   779 => x"e0e2c278",
   780 => x"d4e2c21e",
   781 => x"e2c249bf",
   782 => x"a1c148d4",
   783 => x"ffe27178",
   784 => x"c086c487",
   785 => x"c248ccf7",
   786 => x"cc78e0e2",
   787 => x"ccf7c087",
   788 => x"e0c048bf",
   789 => x"d0f7c080",
   790 => x"dce2c258",
   791 => x"80c148bf",
   792 => x"58e0e2c2",
   793 => x"000dcc27",
   794 => x"bf97bf00",
   795 => x"c2029d4d",
   796 => x"e5c387e5",
   797 => x"dec202ad",
   798 => x"ccf7c087",
   799 => x"a3cb4bbf",
   800 => x"cf4c1149",
   801 => x"d2c105ac",
   802 => x"df497587",
   803 => x"cd89c199",
   804 => x"f0eac291",
   805 => x"4aa3c181",
   806 => x"a3c35112",
   807 => x"c551124a",
   808 => x"51124aa3",
   809 => x"124aa3c7",
   810 => x"4aa3c951",
   811 => x"a3ce5112",
   812 => x"d051124a",
   813 => x"51124aa3",
   814 => x"124aa3d2",
   815 => x"4aa3d451",
   816 => x"a3d65112",
   817 => x"d851124a",
   818 => x"51124aa3",
   819 => x"124aa3dc",
   820 => x"4aa3de51",
   821 => x"7ec15112",
   822 => x"7487fcc0",
   823 => x"0599c849",
   824 => x"7487edc0",
   825 => x"0599d049",
   826 => x"e0c087d3",
   827 => x"ccc00266",
   828 => x"c0497387",
   829 => x"700f66e0",
   830 => x"d3c00298",
   831 => x"c0056e87",
   832 => x"eac287c6",
   833 => x"50c048f0",
   834 => x"bfccf7c0",
   835 => x"87e9c248",
   836 => x"48fdeac2",
   837 => x"c27e50c0",
   838 => x"49bfecea",
   839 => x"bfdce2c2",
   840 => x"04aa714a",
   841 => x"cf87f5fb",
   842 => x"f8ffffff",
   843 => x"d0efc24c",
   844 => x"c8c005bf",
   845 => x"e8eac287",
   846 => x"fac102bf",
   847 => x"d8e2c287",
   848 => x"f9ec49bf",
   849 => x"dce2c287",
   850 => x"48a6c458",
   851 => x"bfd8e2c2",
   852 => x"e8eac278",
   853 => x"dbc002bf",
   854 => x"4966c487",
   855 => x"a9749974",
   856 => x"87c8c002",
   857 => x"c048a6c8",
   858 => x"87e7c078",
   859 => x"c148a6c8",
   860 => x"87dfc078",
   861 => x"cf4966c4",
   862 => x"a999f8ff",
   863 => x"87c8c002",
   864 => x"c048a6cc",
   865 => x"87c5c078",
   866 => x"c148a6cc",
   867 => x"48a6c878",
   868 => x"c87866cc",
   869 => x"dec00566",
   870 => x"4966c487",
   871 => x"eac289c2",
   872 => x"c291bfe0",
   873 => x"48bffcee",
   874 => x"e2c28071",
   875 => x"e2c258d8",
   876 => x"78c048dc",
   877 => x"c087d5f9",
   878 => x"ffffcf48",
   879 => x"f04cf8ff",
   880 => x"264d268e",
   881 => x"264b264c",
   882 => x"0000004f",
   883 => x"00000000",
   884 => x"ffffffff",
   885 => x"00000ddc",
   886 => x"00000de8",
   887 => x"33544146",
   888 => x"20202032",
   889 => x"00000000",
   890 => x"31544146",
   891 => x"20202036",
   892 => x"d4ff1e00",
   893 => x"78ffc348",
   894 => x"4f264868",
   895 => x"48d4ff1e",
   896 => x"ff78ffc3",
   897 => x"e1c048d0",
   898 => x"48d4ff78",
   899 => x"4f2678d4",
   900 => x"48d0ff1e",
   901 => x"2678e0c0",
   902 => x"d4ff1e4f",
   903 => x"99497087",
   904 => x"c087c602",
   905 => x"f105a9fb",
   906 => x"26487187",
   907 => x"5b5e0e4f",
   908 => x"4b710e5c",
   909 => x"f8fe4cc0",
   910 => x"99497087",
   911 => x"87f9c002",
   912 => x"02a9ecc0",
   913 => x"c087f2c0",
   914 => x"c002a9fb",
   915 => x"66cc87eb",
   916 => x"c703acb7",
   917 => x"0266d087",
   918 => x"537187c2",
   919 => x"c2029971",
   920 => x"fe84c187",
   921 => x"497087cb",
   922 => x"87cd0299",
   923 => x"02a9ecc0",
   924 => x"fbc087c7",
   925 => x"d5ff05a9",
   926 => x"0266d087",
   927 => x"97c087c3",
   928 => x"a9ecc07b",
   929 => x"7487c405",
   930 => x"7487c54a",
   931 => x"8a0ac04a",
   932 => x"4c264872",
   933 => x"4f264b26",
   934 => x"87d5fd1e",
   935 => x"f0c04970",
   936 => x"87c904a9",
   937 => x"01a9f9c0",
   938 => x"f0c087c3",
   939 => x"a9c1c189",
   940 => x"c187c904",
   941 => x"c301a9da",
   942 => x"89f7c087",
   943 => x"4f264871",
   944 => x"5c5b5e0e",
   945 => x"86f80e5d",
   946 => x"7ec04c71",
   947 => x"c087edfc",
   948 => x"e0fdc04b",
   949 => x"c049bf97",
   950 => x"87cf04a9",
   951 => x"c187fafc",
   952 => x"e0fdc083",
   953 => x"ab49bf97",
   954 => x"c087f106",
   955 => x"bf97e0fd",
   956 => x"fb87cf02",
   957 => x"497087fb",
   958 => x"87c60299",
   959 => x"05a9ecc0",
   960 => x"4bc087f1",
   961 => x"7087eafb",
   962 => x"87e5fb4d",
   963 => x"fb58a6c8",
   964 => x"4a7087df",
   965 => x"a4c883c1",
   966 => x"49699749",
   967 => x"87da05ad",
   968 => x"9749a4c9",
   969 => x"66c44969",
   970 => x"87ce05a9",
   971 => x"9749a4ca",
   972 => x"05aa4969",
   973 => x"7ec187c4",
   974 => x"ecc087d0",
   975 => x"87c602ad",
   976 => x"05adfbc0",
   977 => x"4bc087c4",
   978 => x"026e7ec1",
   979 => x"fa87f5fe",
   980 => x"487387fe",
   981 => x"4d268ef8",
   982 => x"4b264c26",
   983 => x"00004f26",
   984 => x"1e731e00",
   985 => x"c84bd4ff",
   986 => x"d0ff4a66",
   987 => x"78c5c848",
   988 => x"c148d4ff",
   989 => x"7b1178d4",
   990 => x"f9058ac1",
   991 => x"48d0ff87",
   992 => x"4b2678c4",
   993 => x"5e0e4f26",
   994 => x"0e5d5c5b",
   995 => x"7e7186f8",
   996 => x"efc21e6e",
   997 => x"dce549e0",
   998 => x"7086c487",
   999 => x"e4c40298",
  1000 => x"e8ecc187",
  1001 => x"496e4cbf",
  1002 => x"c887d5fc",
  1003 => x"987058a6",
  1004 => x"c487c505",
  1005 => x"78c148a6",
  1006 => x"c548d0ff",
  1007 => x"48d4ff78",
  1008 => x"c478d5c1",
  1009 => x"89c14966",
  1010 => x"ecc131c6",
  1011 => x"4abf97e0",
  1012 => x"ffb07148",
  1013 => x"ff7808d4",
  1014 => x"78c448d0",
  1015 => x"97dcefc2",
  1016 => x"99d049bf",
  1017 => x"c587dd02",
  1018 => x"48d4ff78",
  1019 => x"c078d6c1",
  1020 => x"48d4ff4a",
  1021 => x"c178ffc3",
  1022 => x"aae0c082",
  1023 => x"ff87f204",
  1024 => x"78c448d0",
  1025 => x"c348d4ff",
  1026 => x"d0ff78ff",
  1027 => x"ff78c548",
  1028 => x"d3c148d4",
  1029 => x"ff78c178",
  1030 => x"78c448d0",
  1031 => x"06acb7c0",
  1032 => x"c287cbc2",
  1033 => x"4bbfe8ef",
  1034 => x"737e748c",
  1035 => x"ddc1029b",
  1036 => x"4dc0c887",
  1037 => x"abb7c08b",
  1038 => x"c887c603",
  1039 => x"c04da3c0",
  1040 => x"dcefc24b",
  1041 => x"d049bf97",
  1042 => x"87cf0299",
  1043 => x"efc21ec0",
  1044 => x"e1e749e0",
  1045 => x"7086c487",
  1046 => x"c287d84c",
  1047 => x"c21ee0e2",
  1048 => x"e749e0ef",
  1049 => x"4c7087d0",
  1050 => x"e2c21e75",
  1051 => x"f0fb49e0",
  1052 => x"7486c887",
  1053 => x"87c5059c",
  1054 => x"cac148c0",
  1055 => x"c21ec187",
  1056 => x"e549e0ef",
  1057 => x"86c487d5",
  1058 => x"fe059b73",
  1059 => x"4c6e87e3",
  1060 => x"06acb7c0",
  1061 => x"efc287d1",
  1062 => x"78c048e0",
  1063 => x"78c080d0",
  1064 => x"efc280f4",
  1065 => x"c078bfec",
  1066 => x"fd01acb7",
  1067 => x"d0ff87f5",
  1068 => x"ff78c548",
  1069 => x"d3c148d4",
  1070 => x"ff78c078",
  1071 => x"78c448d0",
  1072 => x"c2c048c1",
  1073 => x"f848c087",
  1074 => x"264d268e",
  1075 => x"264b264c",
  1076 => x"5b5e0e4f",
  1077 => x"fc0e5d5c",
  1078 => x"c04d7186",
  1079 => x"04ad4c4b",
  1080 => x"c087e8c0",
  1081 => x"741ec0fb",
  1082 => x"87c4029c",
  1083 => x"87c24ac0",
  1084 => x"49724ac1",
  1085 => x"c487dfeb",
  1086 => x"c17e7086",
  1087 => x"c2056e83",
  1088 => x"c14b7587",
  1089 => x"06ab7584",
  1090 => x"6e87d8ff",
  1091 => x"268efc48",
  1092 => x"264c264d",
  1093 => x"0e4f264b",
  1094 => x"0e5c5b5e",
  1095 => x"66cc4b71",
  1096 => x"4c87d802",
  1097 => x"028cf0c0",
  1098 => x"4a7487d8",
  1099 => x"d1028ac1",
  1100 => x"cd028a87",
  1101 => x"c9028a87",
  1102 => x"7387d987",
  1103 => x"87c6f949",
  1104 => x"1e7487d2",
  1105 => x"d9c149c0",
  1106 => x"1e7487ea",
  1107 => x"d9c14973",
  1108 => x"86c887e2",
  1109 => x"4b264c26",
  1110 => x"5e0e4f26",
  1111 => x"0e5d5c5b",
  1112 => x"4c7186fc",
  1113 => x"c291de49",
  1114 => x"714dccf0",
  1115 => x"026d9785",
  1116 => x"c287dcc1",
  1117 => x"49bffcef",
  1118 => x"fd718174",
  1119 => x"7e7087d3",
  1120 => x"c0029848",
  1121 => x"f0c287f2",
  1122 => x"4a704bc0",
  1123 => x"fefe49cb",
  1124 => x"4b7487d2",
  1125 => x"ecc193cc",
  1126 => x"83c483ec",
  1127 => x"7bdcc7c1",
  1128 => x"c4c14974",
  1129 => x"7b7587da",
  1130 => x"97e4ecc1",
  1131 => x"c21e49bf",
  1132 => x"fd49c0f0",
  1133 => x"86c487e1",
  1134 => x"c4c14974",
  1135 => x"49c087c2",
  1136 => x"87ddc5c1",
  1137 => x"48d8efc2",
  1138 => x"c04950c0",
  1139 => x"fc87cce2",
  1140 => x"264d268e",
  1141 => x"264b264c",
  1142 => x"0000004f",
  1143 => x"64616f4c",
  1144 => x"2e676e69",
  1145 => x"1e002e2e",
  1146 => x"4b711e73",
  1147 => x"fcefc249",
  1148 => x"fb7181bf",
  1149 => x"4a7087db",
  1150 => x"87c4029a",
  1151 => x"87dce649",
  1152 => x"48fcefc2",
  1153 => x"497378c0",
  1154 => x"2687fac1",
  1155 => x"1e4f264b",
  1156 => x"4b711e73",
  1157 => x"024aa3c4",
  1158 => x"c187d0c1",
  1159 => x"87dc028a",
  1160 => x"f2c0028a",
  1161 => x"c1058a87",
  1162 => x"efc287d3",
  1163 => x"c102bffc",
  1164 => x"c14887cb",
  1165 => x"c0f0c288",
  1166 => x"87c1c158",
  1167 => x"bffcefc2",
  1168 => x"c289c649",
  1169 => x"c059c0f0",
  1170 => x"c003a9b7",
  1171 => x"efc287ef",
  1172 => x"78c048fc",
  1173 => x"c287e6c0",
  1174 => x"02bff8ef",
  1175 => x"efc287df",
  1176 => x"c148bffc",
  1177 => x"c0f0c280",
  1178 => x"c287d258",
  1179 => x"02bff8ef",
  1180 => x"efc287cb",
  1181 => x"c648bffc",
  1182 => x"c0f0c280",
  1183 => x"c4497358",
  1184 => x"264b2687",
  1185 => x"5b5e0e4f",
  1186 => x"f00e5d5c",
  1187 => x"59a6d086",
  1188 => x"4de0e2c2",
  1189 => x"efc24cc0",
  1190 => x"78c148f8",
  1191 => x"c048a6c8",
  1192 => x"c27e7578",
  1193 => x"48bffcef",
  1194 => x"c106a8c0",
  1195 => x"a6c887c0",
  1196 => x"c27e755c",
  1197 => x"9848e0e2",
  1198 => x"87f2c002",
  1199 => x"c04d66c4",
  1200 => x"cc1ec0fb",
  1201 => x"87c40266",
  1202 => x"87c24cc0",
  1203 => x"49744cc1",
  1204 => x"c487c3e4",
  1205 => x"c17e7086",
  1206 => x"4866c885",
  1207 => x"a6cc80c1",
  1208 => x"fcefc258",
  1209 => x"c503adbf",
  1210 => x"ff056e87",
  1211 => x"4d6e87d1",
  1212 => x"9d754cc0",
  1213 => x"87dcc302",
  1214 => x"1ec0fbc0",
  1215 => x"c70266cc",
  1216 => x"48a6c887",
  1217 => x"87c578c0",
  1218 => x"c148a6c8",
  1219 => x"4966c878",
  1220 => x"c487c3e3",
  1221 => x"487e7086",
  1222 => x"e4c20298",
  1223 => x"81cb4987",
  1224 => x"d0496997",
  1225 => x"d4c10299",
  1226 => x"cc497487",
  1227 => x"ececc191",
  1228 => x"e7c7c181",
  1229 => x"c381c879",
  1230 => x"497451ff",
  1231 => x"f0c291de",
  1232 => x"85714dcc",
  1233 => x"7d97c1c2",
  1234 => x"c049a5c1",
  1235 => x"eac251e0",
  1236 => x"02bf97f0",
  1237 => x"84c187d2",
  1238 => x"c24ba5c2",
  1239 => x"db4af0ea",
  1240 => x"fff6fe49",
  1241 => x"87d9c187",
  1242 => x"c049a5cd",
  1243 => x"c284c151",
  1244 => x"4a6e4ba5",
  1245 => x"f6fe49cb",
  1246 => x"c4c187ea",
  1247 => x"cc497487",
  1248 => x"ececc191",
  1249 => x"dac5c181",
  1250 => x"f0eac279",
  1251 => x"d802bf97",
  1252 => x"de497487",
  1253 => x"c284c191",
  1254 => x"714bccf0",
  1255 => x"f0eac283",
  1256 => x"fe49dd4a",
  1257 => x"d887fdf5",
  1258 => x"de4b7487",
  1259 => x"ccf0c293",
  1260 => x"49a3cb83",
  1261 => x"84c151c0",
  1262 => x"cb4a6e73",
  1263 => x"e3f5fe49",
  1264 => x"4866c887",
  1265 => x"a6cc80c1",
  1266 => x"03acc758",
  1267 => x"6e87c5c0",
  1268 => x"87e4fc05",
  1269 => x"c003acc7",
  1270 => x"efc287e4",
  1271 => x"78c048f8",
  1272 => x"91cc4974",
  1273 => x"81ececc1",
  1274 => x"79dac5c1",
  1275 => x"91de4974",
  1276 => x"81ccf0c2",
  1277 => x"84c151c0",
  1278 => x"ff04acc7",
  1279 => x"eec187dc",
  1280 => x"50c048c8",
  1281 => x"d1c180f7",
  1282 => x"d0c140f5",
  1283 => x"80c878e8",
  1284 => x"78cfc8c1",
  1285 => x"c04966cc",
  1286 => x"f087e5fa",
  1287 => x"264d268e",
  1288 => x"264b264c",
  1289 => x"0000004f",
  1290 => x"61422080",
  1291 => x"1e006b63",
  1292 => x"4b711e73",
  1293 => x"c191cc49",
  1294 => x"c881ecec",
  1295 => x"ecc14aa1",
  1296 => x"501248e0",
  1297 => x"c04aa1c9",
  1298 => x"1248e0fd",
  1299 => x"c181ca50",
  1300 => x"1148e4ec",
  1301 => x"e4ecc150",
  1302 => x"1e49bf97",
  1303 => x"f6f249c0",
  1304 => x"f8497387",
  1305 => x"8efc87df",
  1306 => x"4f264b26",
  1307 => x"c049c01e",
  1308 => x"2687eefa",
  1309 => x"4a711e4f",
  1310 => x"c191cc49",
  1311 => x"c881ecec",
  1312 => x"d8efc281",
  1313 => x"c0501148",
  1314 => x"fe49a2f0",
  1315 => x"c087fdef",
  1316 => x"87c7d749",
  1317 => x"ff1e4f26",
  1318 => x"ffc34ad4",
  1319 => x"48d0ff7a",
  1320 => x"de78e1c0",
  1321 => x"487a717a",
  1322 => x"7028b7c8",
  1323 => x"d048717a",
  1324 => x"7a7028b7",
  1325 => x"b7d84871",
  1326 => x"ff7a7028",
  1327 => x"e0c048d0",
  1328 => x"0e4f2678",
  1329 => x"5d5c5b5e",
  1330 => x"7186f40e",
  1331 => x"91cc494d",
  1332 => x"81ececc1",
  1333 => x"ca4aa1c8",
  1334 => x"a6c47ea1",
  1335 => x"d4efc248",
  1336 => x"976e78bf",
  1337 => x"66c44bbf",
  1338 => x"122c734c",
  1339 => x"58a6cc48",
  1340 => x"84c19c70",
  1341 => x"699781c9",
  1342 => x"04acb749",
  1343 => x"4cc087c2",
  1344 => x"4abf976e",
  1345 => x"724966c8",
  1346 => x"c4b9ff31",
  1347 => x"48749966",
  1348 => x"4a703072",
  1349 => x"d8efc2b1",
  1350 => x"f9fd7159",
  1351 => x"c21ec787",
  1352 => x"1ebff4ef",
  1353 => x"1eececc1",
  1354 => x"97d8efc2",
  1355 => x"f4c149bf",
  1356 => x"c0497587",
  1357 => x"e887c9f6",
  1358 => x"264d268e",
  1359 => x"264b264c",
  1360 => x"1e731e4f",
  1361 => x"fd494b71",
  1362 => x"497387f9",
  1363 => x"2687f4fd",
  1364 => x"1e4f264b",
  1365 => x"4b711e73",
  1366 => x"024aa3c2",
  1367 => x"8ac187d6",
  1368 => x"87e2c005",
  1369 => x"bff4efc2",
  1370 => x"4887db02",
  1371 => x"efc288c1",
  1372 => x"87d258f8",
  1373 => x"bff8efc2",
  1374 => x"c287cb02",
  1375 => x"48bff4ef",
  1376 => x"efc280c1",
  1377 => x"1ec758f8",
  1378 => x"bff4efc2",
  1379 => x"ececc11e",
  1380 => x"d8efc21e",
  1381 => x"cc49bf97",
  1382 => x"c0497387",
  1383 => x"f487e1f4",
  1384 => x"264b268e",
  1385 => x"5b5e0e4f",
  1386 => x"ff0e5d5c",
  1387 => x"e4c086cc",
  1388 => x"a6cc59a6",
  1389 => x"c478c048",
  1390 => x"c478c080",
  1391 => x"66c8c180",
  1392 => x"c180c478",
  1393 => x"c180c478",
  1394 => x"f8efc278",
  1395 => x"e078c148",
  1396 => x"c4e187ea",
  1397 => x"87d9e087",
  1398 => x"fbc04c70",
  1399 => x"f3c102ac",
  1400 => x"66e0c087",
  1401 => x"87e8c105",
  1402 => x"4a66c4c1",
  1403 => x"7e6a82c4",
  1404 => x"48fce8c1",
  1405 => x"4120496e",
  1406 => x"51104120",
  1407 => x"4866c4c1",
  1408 => x"78efd0c1",
  1409 => x"81c7496a",
  1410 => x"c4c15174",
  1411 => x"81c84966",
  1412 => x"a6d851c1",
  1413 => x"c178c248",
  1414 => x"c94966c4",
  1415 => x"c151c081",
  1416 => x"ca4966c4",
  1417 => x"c151c081",
  1418 => x"6a1ed81e",
  1419 => x"ff81c849",
  1420 => x"c887fadf",
  1421 => x"66c8c186",
  1422 => x"01a8c048",
  1423 => x"a6d087c7",
  1424 => x"cf78c148",
  1425 => x"66c8c187",
  1426 => x"d888c148",
  1427 => x"87c458a6",
  1428 => x"87c5dfff",
  1429 => x"cd029c74",
  1430 => x"66d087d9",
  1431 => x"66ccc148",
  1432 => x"cecd03a8",
  1433 => x"48a6c887",
  1434 => x"ff7e78c0",
  1435 => x"7087c2de",
  1436 => x"acd0c14c",
  1437 => x"87e7c205",
  1438 => x"6e48a6c4",
  1439 => x"87d8e078",
  1440 => x"cc487e70",
  1441 => x"c506a866",
  1442 => x"48a6cc87",
  1443 => x"ddff786e",
  1444 => x"4c7087df",
  1445 => x"05acecc0",
  1446 => x"d087eec1",
  1447 => x"91cc4966",
  1448 => x"8166c4c1",
  1449 => x"6a4aa1c4",
  1450 => x"4aa1c84d",
  1451 => x"d1c1526e",
  1452 => x"dcff79f5",
  1453 => x"4c7087fb",
  1454 => x"87d9029c",
  1455 => x"02acfbc0",
  1456 => x"557487d3",
  1457 => x"87e9dcff",
  1458 => x"029c4c70",
  1459 => x"fbc087c7",
  1460 => x"edff05ac",
  1461 => x"55e0c087",
  1462 => x"c055c1c2",
  1463 => x"e0c07d97",
  1464 => x"66c44866",
  1465 => x"87db05a8",
  1466 => x"d44866d0",
  1467 => x"ca04a866",
  1468 => x"4866d087",
  1469 => x"a6d480c1",
  1470 => x"d487c858",
  1471 => x"88c14866",
  1472 => x"ff58a6d8",
  1473 => x"7087eadb",
  1474 => x"acd0c14c",
  1475 => x"dc87c905",
  1476 => x"80c14866",
  1477 => x"58a6e0c0",
  1478 => x"02acd0c1",
  1479 => x"6e87d9fd",
  1480 => x"66e0c048",
  1481 => x"eac905a8",
  1482 => x"a6e4c087",
  1483 => x"7478c048",
  1484 => x"88fbc048",
  1485 => x"7058a6c8",
  1486 => x"dcc90298",
  1487 => x"88cb4887",
  1488 => x"7058a6c8",
  1489 => x"cec10298",
  1490 => x"88c94887",
  1491 => x"7058a6c8",
  1492 => x"fec30298",
  1493 => x"88c44887",
  1494 => x"7058a6c8",
  1495 => x"87cf0298",
  1496 => x"c888c148",
  1497 => x"987058a6",
  1498 => x"87e7c302",
  1499 => x"c887dbc8",
  1500 => x"f0c048a6",
  1501 => x"f8d9ff78",
  1502 => x"c04c7087",
  1503 => x"c302acec",
  1504 => x"5ca6cc87",
  1505 => x"02acecc0",
  1506 => x"d9ff87cd",
  1507 => x"4c7087e3",
  1508 => x"05acecc0",
  1509 => x"c087f3ff",
  1510 => x"c002acec",
  1511 => x"d9ff87c4",
  1512 => x"1ec087cf",
  1513 => x"66d81eca",
  1514 => x"c191cc49",
  1515 => x"714866cc",
  1516 => x"58a6cc80",
  1517 => x"c44866c8",
  1518 => x"58a6d080",
  1519 => x"49bf66cc",
  1520 => x"87e9d9ff",
  1521 => x"1ede1ec1",
  1522 => x"49bf66d4",
  1523 => x"87ddd9ff",
  1524 => x"497086d0",
  1525 => x"8808c048",
  1526 => x"58a6ecc0",
  1527 => x"c006a8c0",
  1528 => x"e8c087ee",
  1529 => x"a8dd4866",
  1530 => x"87e4c003",
  1531 => x"49bf66c4",
  1532 => x"8166e8c0",
  1533 => x"c051e0c0",
  1534 => x"c14966e8",
  1535 => x"bf66c481",
  1536 => x"51c1c281",
  1537 => x"4966e8c0",
  1538 => x"66c481c2",
  1539 => x"51c081bf",
  1540 => x"d0c1486e",
  1541 => x"496e78ef",
  1542 => x"66d881c8",
  1543 => x"c9496e51",
  1544 => x"5166dc81",
  1545 => x"81ca496e",
  1546 => x"d85166c8",
  1547 => x"80c14866",
  1548 => x"d058a6dc",
  1549 => x"66d44866",
  1550 => x"cbc004a8",
  1551 => x"4866d087",
  1552 => x"a6d480c1",
  1553 => x"87d1c558",
  1554 => x"c14866d4",
  1555 => x"58a6d888",
  1556 => x"ff87c6c5",
  1557 => x"c087c1d9",
  1558 => x"ff58a6ec",
  1559 => x"c087f9d8",
  1560 => x"c058a6f0",
  1561 => x"c005a8ec",
  1562 => x"48a687c9",
  1563 => x"7866e8c0",
  1564 => x"ff87c4c0",
  1565 => x"d087fad5",
  1566 => x"91cc4966",
  1567 => x"4866c4c1",
  1568 => x"a6c88071",
  1569 => x"4a66c458",
  1570 => x"66c482c8",
  1571 => x"c081ca49",
  1572 => x"c05166e8",
  1573 => x"c14966ec",
  1574 => x"66e8c081",
  1575 => x"7148c189",
  1576 => x"c1497030",
  1577 => x"7a977189",
  1578 => x"bfd4efc2",
  1579 => x"66e8c049",
  1580 => x"4a6a9729",
  1581 => x"c0987148",
  1582 => x"c458a6f4",
  1583 => x"80c44866",
  1584 => x"c858a6cc",
  1585 => x"c04dbf66",
  1586 => x"6e4866e0",
  1587 => x"c5c002a8",
  1588 => x"c07ec087",
  1589 => x"7ec187c2",
  1590 => x"e0c01e6e",
  1591 => x"ff49751e",
  1592 => x"c887cad5",
  1593 => x"c04c7086",
  1594 => x"c106acb7",
  1595 => x"857487d4",
  1596 => x"49bf66c8",
  1597 => x"7581e0c0",
  1598 => x"e9c14b89",
  1599 => x"fe714ac8",
  1600 => x"c287e1e0",
  1601 => x"c07e7585",
  1602 => x"c14866e4",
  1603 => x"a6e8c080",
  1604 => x"66f0c058",
  1605 => x"7081c149",
  1606 => x"c5c002a9",
  1607 => x"c04dc087",
  1608 => x"4dc187c2",
  1609 => x"66cc1e75",
  1610 => x"e0c049bf",
  1611 => x"8966c481",
  1612 => x"66c81e71",
  1613 => x"f4d3ff49",
  1614 => x"c086c887",
  1615 => x"ff01a8b7",
  1616 => x"e4c087c5",
  1617 => x"d3c00266",
  1618 => x"4966c487",
  1619 => x"e4c081c9",
  1620 => x"66c45166",
  1621 => x"c3d3c148",
  1622 => x"87cec078",
  1623 => x"c94966c4",
  1624 => x"c451c281",
  1625 => x"d5c14866",
  1626 => x"66d078c1",
  1627 => x"a866d448",
  1628 => x"87cbc004",
  1629 => x"c14866d0",
  1630 => x"58a6d480",
  1631 => x"d487dac0",
  1632 => x"88c14866",
  1633 => x"c058a6d8",
  1634 => x"d2ff87cf",
  1635 => x"4c7087cb",
  1636 => x"ff87c6c0",
  1637 => x"7087c2d2",
  1638 => x"4866dc4c",
  1639 => x"e0c080c1",
  1640 => x"9c7458a6",
  1641 => x"87cbc002",
  1642 => x"c14866d0",
  1643 => x"04a866cc",
  1644 => x"d087f2f2",
  1645 => x"a8c74866",
  1646 => x"87e1c003",
  1647 => x"c24c66d0",
  1648 => x"c048f8ef",
  1649 => x"cc497478",
  1650 => x"66c4c191",
  1651 => x"4aa1c481",
  1652 => x"52c04a6a",
  1653 => x"c784c179",
  1654 => x"e2ff04ac",
  1655 => x"66e0c087",
  1656 => x"87e2c002",
  1657 => x"4966c4c1",
  1658 => x"c181d4c1",
  1659 => x"c14a66c4",
  1660 => x"52c082dc",
  1661 => x"79f5d1c1",
  1662 => x"4966c4c1",
  1663 => x"c181d8c1",
  1664 => x"c079cce9",
  1665 => x"c4c187d6",
  1666 => x"d4c14966",
  1667 => x"66c4c181",
  1668 => x"82d8c14a",
  1669 => x"7ad4e9c1",
  1670 => x"79ecd1c1",
  1671 => x"4966c4c1",
  1672 => x"c181e0c1",
  1673 => x"ff79d3d5",
  1674 => x"cc87e5cf",
  1675 => x"ccff4866",
  1676 => x"264d268e",
  1677 => x"264b264c",
  1678 => x"0000004f",
  1679 => x"64616f4c",
  1680 => x"202e2a20",
  1681 => x"00000000",
  1682 => x"0000203a",
  1683 => x"61422080",
  1684 => x"00006b63",
  1685 => x"78452080",
  1686 => x"1e007469",
  1687 => x"efc21ec7",
  1688 => x"c11ebff4",
  1689 => x"c21eecec",
  1690 => x"bf97d8ef",
  1691 => x"87f5ec49",
  1692 => x"49ececc1",
  1693 => x"87d6e2c0",
  1694 => x"4f268ef4",
  1695 => x"c81e731e",
  1696 => x"eec187c3",
  1697 => x"ecc148c4",
  1698 => x"e8fe78cc",
  1699 => x"e1c049a0",
  1700 => x"49c787fc",
  1701 => x"87e8e0c0",
  1702 => x"e2c049c1",
  1703 => x"d4ff87c3",
  1704 => x"78ffc348",
  1705 => x"48c0f0c2",
  1706 => x"e3fe50c0",
  1707 => x"987087de",
  1708 => x"fe87cd02",
  1709 => x"7087daed",
  1710 => x"87c40298",
  1711 => x"87c24ac1",
  1712 => x"9a724ac0",
  1713 => x"c187c802",
  1714 => x"fe49d8ec",
  1715 => x"c287d8d7",
  1716 => x"c048f4ef",
  1717 => x"d8efc278",
  1718 => x"4950c048",
  1719 => x"c087fcfd",
  1720 => x"7087d5f5",
  1721 => x"cb029b4b",
  1722 => x"c8eec187",
  1723 => x"df49c75b",
  1724 => x"87c687ce",
  1725 => x"e0c049c0",
  1726 => x"c2c387e7",
  1727 => x"c8e2c087",
  1728 => x"dcefc087",
  1729 => x"87f5ff87",
  1730 => x"4f264b26",
  1731 => x"746f6f42",
  1732 => x"2e676e69",
  1733 => x"00002e2e",
  1734 => x"4f204453",
  1735 => x"0000004b",
  1736 => x"00000000",
  1737 => x"00000000",
  1738 => x"00000001",
  1739 => x"0000115a",
  1740 => x"00002c0c",
  1741 => x"00000000",
  1742 => x"0000115a",
  1743 => x"00002c2a",
  1744 => x"00000000",
  1745 => x"0000115a",
  1746 => x"00002c48",
  1747 => x"00000000",
  1748 => x"0000115a",
  1749 => x"00002c66",
  1750 => x"00000000",
  1751 => x"0000115a",
  1752 => x"00002c84",
  1753 => x"00000000",
  1754 => x"0000115a",
  1755 => x"00002ca2",
  1756 => x"00000000",
  1757 => x"0000115a",
  1758 => x"00002cc0",
  1759 => x"00000000",
  1760 => x"00001475",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"0000120f",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"db86fc1e",
  1767 => x"fc7e7087",
  1768 => x"1e4f268e",
  1769 => x"c048f0fe",
  1770 => x"7909cd78",
  1771 => x"1e4f2609",
  1772 => x"49d8eec1",
  1773 => x"4f2687ed",
  1774 => x"bff0fe1e",
  1775 => x"1e4f2648",
  1776 => x"c148f0fe",
  1777 => x"1e4f2678",
  1778 => x"c048f0fe",
  1779 => x"1e4f2678",
  1780 => x"52c04a71",
  1781 => x"0e4f2651",
  1782 => x"5d5c5b5e",
  1783 => x"7186f40e",
  1784 => x"7e6d974d",
  1785 => x"974ca5c1",
  1786 => x"a6c8486c",
  1787 => x"c4486e58",
  1788 => x"c505a866",
  1789 => x"c048ff87",
  1790 => x"caff87e6",
  1791 => x"49a5c287",
  1792 => x"714b6c97",
  1793 => x"6b974ba3",
  1794 => x"7e6c974b",
  1795 => x"80c1486e",
  1796 => x"c758a6c8",
  1797 => x"58a6cc98",
  1798 => x"fe7c9770",
  1799 => x"487387e1",
  1800 => x"4d268ef4",
  1801 => x"4b264c26",
  1802 => x"5e0e4f26",
  1803 => x"f40e5c5b",
  1804 => x"d84c7186",
  1805 => x"ffc34a66",
  1806 => x"4ba4c29a",
  1807 => x"73496c97",
  1808 => x"517249a1",
  1809 => x"6e7e6c97",
  1810 => x"c880c148",
  1811 => x"98c758a6",
  1812 => x"7058a6cc",
  1813 => x"268ef454",
  1814 => x"264b264c",
  1815 => x"86fc1e4f",
  1816 => x"e087e4fd",
  1817 => x"c0494abf",
  1818 => x"0299c0e0",
  1819 => x"1e7287cb",
  1820 => x"49e0f3c2",
  1821 => x"c487f3fe",
  1822 => x"87fcfc86",
  1823 => x"fefc7e70",
  1824 => x"268efc87",
  1825 => x"f3c21e4f",
  1826 => x"c2fd49e0",
  1827 => x"ddf1c187",
  1828 => x"87cffc49",
  1829 => x"2687edc3",
  1830 => x"5b5e0e4f",
  1831 => x"fc0e5d5c",
  1832 => x"ff7e7186",
  1833 => x"f3c24dd4",
  1834 => x"eafc49e0",
  1835 => x"c04b7087",
  1836 => x"c204abb7",
  1837 => x"f0c387f8",
  1838 => x"87c905ab",
  1839 => x"48fcf5c1",
  1840 => x"d9c278c1",
  1841 => x"abe0c387",
  1842 => x"c187c905",
  1843 => x"c148c0f6",
  1844 => x"87cac278",
  1845 => x"bfc0f6c1",
  1846 => x"c287c602",
  1847 => x"c24ca3c0",
  1848 => x"c14c7387",
  1849 => x"02bffcf5",
  1850 => x"7487e0c0",
  1851 => x"29b7c449",
  1852 => x"d8f7c191",
  1853 => x"cf4a7481",
  1854 => x"c192c29a",
  1855 => x"70307248",
  1856 => x"72baff4a",
  1857 => x"70986948",
  1858 => x"7487db79",
  1859 => x"29b7c449",
  1860 => x"d8f7c191",
  1861 => x"cf4a7481",
  1862 => x"c392c29a",
  1863 => x"70307248",
  1864 => x"b069484a",
  1865 => x"056e7970",
  1866 => x"ff87e7c0",
  1867 => x"e1c848d0",
  1868 => x"c17dc578",
  1869 => x"02bfc0f6",
  1870 => x"e0c387c3",
  1871 => x"fcf5c17d",
  1872 => x"87c302bf",
  1873 => x"737df0c3",
  1874 => x"48d0ff7d",
  1875 => x"c078e1c8",
  1876 => x"f6c178e0",
  1877 => x"78c048c0",
  1878 => x"48fcf5c1",
  1879 => x"f3c278c0",
  1880 => x"f2f949e0",
  1881 => x"c04b7087",
  1882 => x"fd03abb7",
  1883 => x"48c087c8",
  1884 => x"4d268efc",
  1885 => x"4b264c26",
  1886 => x"00004f26",
  1887 => x"00000000",
  1888 => x"00000000",
  1889 => x"724ac01e",
  1890 => x"c191c449",
  1891 => x"c081d8f7",
  1892 => x"d082c179",
  1893 => x"ee04aab7",
  1894 => x"0e4f2687",
  1895 => x"5d5c5b5e",
  1896 => x"f84d710e",
  1897 => x"4a7587e1",
  1898 => x"922ab7c4",
  1899 => x"82d8f7c1",
  1900 => x"9ccf4c75",
  1901 => x"496a94c2",
  1902 => x"c32b744b",
  1903 => x"7448c29b",
  1904 => x"ff4c7030",
  1905 => x"714874bc",
  1906 => x"f77a7098",
  1907 => x"487387f1",
  1908 => x"4c264d26",
  1909 => x"4f264b26",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"00000000",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"00000000",
  1926 => x"48d0ff1e",
  1927 => x"7178e1c8",
  1928 => x"08d4ff48",
  1929 => x"1e4f2678",
  1930 => x"c848d0ff",
  1931 => x"487178e1",
  1932 => x"7808d4ff",
  1933 => x"ff4866c4",
  1934 => x"267808d4",
  1935 => x"4a711e4f",
  1936 => x"1e4966c4",
  1937 => x"deff4972",
  1938 => x"48d0ff87",
  1939 => x"fc78e0c0",
  1940 => x"1e4f268e",
  1941 => x"4b711e73",
  1942 => x"1e4966c8",
  1943 => x"e0c14a73",
  1944 => x"d8ff49a2",
  1945 => x"268efc87",
  1946 => x"1e4f264b",
  1947 => x"c848d0ff",
  1948 => x"487178c9",
  1949 => x"7808d4ff",
  1950 => x"711e4f26",
  1951 => x"87eb494a",
  1952 => x"c848d0ff",
  1953 => x"1e4f2678",
  1954 => x"4b711e73",
  1955 => x"bff8f3c2",
  1956 => x"c287c302",
  1957 => x"d0ff87eb",
  1958 => x"78c9c848",
  1959 => x"e0c04873",
  1960 => x"08d4ffb0",
  1961 => x"ecf3c278",
  1962 => x"c878c048",
  1963 => x"87c50266",
  1964 => x"c249ffc3",
  1965 => x"c249c087",
  1966 => x"cc59f4f3",
  1967 => x"87c60266",
  1968 => x"4ad5d5c5",
  1969 => x"ffcf87c4",
  1970 => x"f3c24aff",
  1971 => x"f3c25af8",
  1972 => x"78c148f8",
  1973 => x"4f264b26",
  1974 => x"5c5b5e0e",
  1975 => x"4d710e5d",
  1976 => x"bff4f3c2",
  1977 => x"029d754b",
  1978 => x"c84987cb",
  1979 => x"c0fac191",
  1980 => x"c482714a",
  1981 => x"c0fec187",
  1982 => x"124cc04a",
  1983 => x"c2997349",
  1984 => x"48bff0f3",
  1985 => x"d4ffb871",
  1986 => x"b7c17808",
  1987 => x"b7c8842b",
  1988 => x"87e704ac",
  1989 => x"bfecf3c2",
  1990 => x"c280c848",
  1991 => x"2658f0f3",
  1992 => x"264c264d",
  1993 => x"1e4f264b",
  1994 => x"4b711e73",
  1995 => x"029a4a13",
  1996 => x"497287cb",
  1997 => x"1387e1fe",
  1998 => x"f5059a4a",
  1999 => x"264b2687",
  2000 => x"f3c21e4f",
  2001 => x"c249bfec",
  2002 => x"c148ecf3",
  2003 => x"c0c478a1",
  2004 => x"db03a9b7",
  2005 => x"48d4ff87",
  2006 => x"bff0f3c2",
  2007 => x"ecf3c278",
  2008 => x"f3c249bf",
  2009 => x"a1c148ec",
  2010 => x"b7c0c478",
  2011 => x"87e504a9",
  2012 => x"c848d0ff",
  2013 => x"f8f3c278",
  2014 => x"2678c048",
  2015 => x"0000004f",
  2016 => x"00000000",
  2017 => x"00000000",
  2018 => x"5f000000",
  2019 => x"0000005f",
  2020 => x"00030300",
  2021 => x"00000303",
  2022 => x"147f7f14",
  2023 => x"00147f7f",
  2024 => x"6b2e2400",
  2025 => x"00123a6b",
  2026 => x"18366a4c",
  2027 => x"0032566c",
  2028 => x"594f7e30",
  2029 => x"40683a77",
  2030 => x"07040000",
  2031 => x"00000003",
  2032 => x"3e1c0000",
  2033 => x"00004163",
  2034 => x"63410000",
  2035 => x"00001c3e",
  2036 => x"1c3e2a08",
  2037 => x"082a3e1c",
  2038 => x"3e080800",
  2039 => x"0008083e",
  2040 => x"e0800000",
  2041 => x"00000060",
  2042 => x"08080800",
  2043 => x"00080808",
  2044 => x"60000000",
  2045 => x"00000060",
  2046 => x"18306040",
  2047 => x"0103060c",
  2048 => x"597f3e00",
  2049 => x"003e7f4d",
  2050 => x"7f060400",
  2051 => x"0000007f",
  2052 => x"71634200",
  2053 => x"00464f59",
  2054 => x"49632200",
  2055 => x"00367f49",
  2056 => x"13161c18",
  2057 => x"00107f7f",
  2058 => x"45672700",
  2059 => x"00397d45",
  2060 => x"4b7e3c00",
  2061 => x"00307949",
  2062 => x"71010100",
  2063 => x"00070f79",
  2064 => x"497f3600",
  2065 => x"00367f49",
  2066 => x"494f0600",
  2067 => x"001e3f69",
  2068 => x"66000000",
  2069 => x"00000066",
  2070 => x"e6800000",
  2071 => x"00000066",
  2072 => x"14080800",
  2073 => x"00222214",
  2074 => x"14141400",
  2075 => x"00141414",
  2076 => x"14222200",
  2077 => x"00080814",
  2078 => x"51030200",
  2079 => x"00060f59",
  2080 => x"5d417f3e",
  2081 => x"001e1f55",
  2082 => x"097f7e00",
  2083 => x"007e7f09",
  2084 => x"497f7f00",
  2085 => x"00367f49",
  2086 => x"633e1c00",
  2087 => x"00414141",
  2088 => x"417f7f00",
  2089 => x"001c3e63",
  2090 => x"497f7f00",
  2091 => x"00414149",
  2092 => x"097f7f00",
  2093 => x"00010109",
  2094 => x"417f3e00",
  2095 => x"007a7b49",
  2096 => x"087f7f00",
  2097 => x"007f7f08",
  2098 => x"7f410000",
  2099 => x"0000417f",
  2100 => x"40602000",
  2101 => x"003f7f40",
  2102 => x"1c087f7f",
  2103 => x"00416336",
  2104 => x"407f7f00",
  2105 => x"00404040",
  2106 => x"0c067f7f",
  2107 => x"007f7f06",
  2108 => x"0c067f7f",
  2109 => x"007f7f18",
  2110 => x"417f3e00",
  2111 => x"003e7f41",
  2112 => x"097f7f00",
  2113 => x"00060f09",
  2114 => x"61417f3e",
  2115 => x"00407e7f",
  2116 => x"097f7f00",
  2117 => x"00667f19",
  2118 => x"4d6f2600",
  2119 => x"00327b59",
  2120 => x"7f010100",
  2121 => x"0001017f",
  2122 => x"407f3f00",
  2123 => x"003f7f40",
  2124 => x"703f0f00",
  2125 => x"000f3f70",
  2126 => x"18307f7f",
  2127 => x"007f7f30",
  2128 => x"1c366341",
  2129 => x"4163361c",
  2130 => x"7c060301",
  2131 => x"0103067c",
  2132 => x"4d597161",
  2133 => x"00414347",
  2134 => x"7f7f0000",
  2135 => x"00004141",
  2136 => x"0c060301",
  2137 => x"40603018",
  2138 => x"41410000",
  2139 => x"00007f7f",
  2140 => x"03060c08",
  2141 => x"00080c06",
  2142 => x"80808080",
  2143 => x"00808080",
  2144 => x"03000000",
  2145 => x"00000407",
  2146 => x"54742000",
  2147 => x"00787c54",
  2148 => x"447f7f00",
  2149 => x"00387c44",
  2150 => x"447c3800",
  2151 => x"00004444",
  2152 => x"447c3800",
  2153 => x"007f7f44",
  2154 => x"547c3800",
  2155 => x"00185c54",
  2156 => x"7f7e0400",
  2157 => x"00000505",
  2158 => x"a4bc1800",
  2159 => x"007cfca4",
  2160 => x"047f7f00",
  2161 => x"00787c04",
  2162 => x"3d000000",
  2163 => x"0000407d",
  2164 => x"80808000",
  2165 => x"00007dfd",
  2166 => x"107f7f00",
  2167 => x"00446c38",
  2168 => x"3f000000",
  2169 => x"0000407f",
  2170 => x"180c7c7c",
  2171 => x"00787c0c",
  2172 => x"047c7c00",
  2173 => x"00787c04",
  2174 => x"447c3800",
  2175 => x"00387c44",
  2176 => x"24fcfc00",
  2177 => x"00183c24",
  2178 => x"243c1800",
  2179 => x"00fcfc24",
  2180 => x"047c7c00",
  2181 => x"00080c04",
  2182 => x"545c4800",
  2183 => x"00207454",
  2184 => x"7f3f0400",
  2185 => x"00004444",
  2186 => x"407c3c00",
  2187 => x"007c7c40",
  2188 => x"603c1c00",
  2189 => x"001c3c60",
  2190 => x"30607c3c",
  2191 => x"003c7c60",
  2192 => x"10386c44",
  2193 => x"00446c38",
  2194 => x"e0bc1c00",
  2195 => x"001c3c60",
  2196 => x"74644400",
  2197 => x"00444c5c",
  2198 => x"3e080800",
  2199 => x"00414177",
  2200 => x"7f000000",
  2201 => x"0000007f",
  2202 => x"77414100",
  2203 => x"0008083e",
  2204 => x"03010102",
  2205 => x"00010202",
  2206 => x"7f7f7f7f",
  2207 => x"007f7f7f",
  2208 => x"1c1c0808",
  2209 => x"7f7f3e3e",
  2210 => x"3e3e7f7f",
  2211 => x"08081c1c",
  2212 => x"7c181000",
  2213 => x"0010187c",
  2214 => x"7c301000",
  2215 => x"0010307c",
  2216 => x"60603010",
  2217 => x"00061e78",
  2218 => x"183c6642",
  2219 => x"0042663c",
  2220 => x"c26a3878",
  2221 => x"00386cc6",
  2222 => x"60000060",
  2223 => x"00600000",
  2224 => x"5c5b5e0e",
  2225 => x"86fc0e5d",
  2226 => x"f4c27e71",
  2227 => x"c04cbfc0",
  2228 => x"c41ec04b",
  2229 => x"c402ab66",
  2230 => x"c24dc087",
  2231 => x"754dc187",
  2232 => x"ee49731e",
  2233 => x"86c887e1",
  2234 => x"ef49e0c0",
  2235 => x"a4c487ea",
  2236 => x"f0496a4a",
  2237 => x"c8f187f1",
  2238 => x"c184cc87",
  2239 => x"abb7c883",
  2240 => x"87cdff04",
  2241 => x"4d268efc",
  2242 => x"4b264c26",
  2243 => x"711e4f26",
  2244 => x"c4f4c24a",
  2245 => x"c4f4c25a",
  2246 => x"4978c748",
  2247 => x"2687e1fe",
  2248 => x"1e731e4f",
  2249 => x"b7c04a71",
  2250 => x"87d303aa",
  2251 => x"bfc4d9c2",
  2252 => x"c187c405",
  2253 => x"c087c24b",
  2254 => x"c8d9c24b",
  2255 => x"c287c45b",
  2256 => x"fc5ac8d9",
  2257 => x"c4d9c248",
  2258 => x"c14a78bf",
  2259 => x"a2c0c19a",
  2260 => x"87e6ec49",
  2261 => x"4f264b26",
  2262 => x"c44a711e",
  2263 => x"49721e66",
  2264 => x"fc87f0eb",
  2265 => x"1e4f268e",
  2266 => x"c348d4ff",
  2267 => x"d0ff78ff",
  2268 => x"78e1c048",
  2269 => x"c148d4ff",
  2270 => x"c4487178",
  2271 => x"08d4ff30",
  2272 => x"48d0ff78",
  2273 => x"2678e0c0",
  2274 => x"5b5e0e4f",
  2275 => x"f00e5d5c",
  2276 => x"48a6c886",
  2277 => x"ec4d78c0",
  2278 => x"80fc7ebf",
  2279 => x"bfc0f4c2",
  2280 => x"4cbfe878",
  2281 => x"bfc4d9c2",
  2282 => x"87ede349",
  2283 => x"ca49eecb",
  2284 => x"4b7087d6",
  2285 => x"e2e749c7",
  2286 => x"05987087",
  2287 => x"496e87c8",
  2288 => x"c10299c1",
  2289 => x"4dc187c1",
  2290 => x"c27ebfec",
  2291 => x"49bfc4d9",
  2292 => x"7387c6e3",
  2293 => x"87fcc949",
  2294 => x"d7029870",
  2295 => x"fcd8c287",
  2296 => x"b9c149bf",
  2297 => x"59c0d9c2",
  2298 => x"87fbfd71",
  2299 => x"c949eecb",
  2300 => x"4b7087d6",
  2301 => x"e2e649c7",
  2302 => x"05987087",
  2303 => x"6e87c7ff",
  2304 => x"0599c149",
  2305 => x"7587fffe",
  2306 => x"e3c0029d",
  2307 => x"c4d9c287",
  2308 => x"bac14abf",
  2309 => x"5ac8d9c2",
  2310 => x"0a7a0afc",
  2311 => x"c0c19ac1",
  2312 => x"d5e949a2",
  2313 => x"49dac187",
  2314 => x"c887f0e5",
  2315 => x"78c148a6",
  2316 => x"bfc4d9c2",
  2317 => x"87e9c005",
  2318 => x"ffc34974",
  2319 => x"c01e7199",
  2320 => x"87d4fc49",
  2321 => x"b7c84974",
  2322 => x"c11e7129",
  2323 => x"87c8fc49",
  2324 => x"fdc386c8",
  2325 => x"87c3e549",
  2326 => x"e449fac3",
  2327 => x"d1c787fd",
  2328 => x"c3497487",
  2329 => x"b7c899ff",
  2330 => x"74b4712c",
  2331 => x"87df029c",
  2332 => x"bfc0d9c2",
  2333 => x"87dcc749",
  2334 => x"c0059870",
  2335 => x"4cc087c4",
  2336 => x"e0c287d3",
  2337 => x"87c0c749",
  2338 => x"58c4d9c2",
  2339 => x"c287c6c0",
  2340 => x"c048c0d9",
  2341 => x"c8497478",
  2342 => x"87ce0599",
  2343 => x"e349f5c3",
  2344 => x"497087f9",
  2345 => x"c00299c2",
  2346 => x"f4c287e9",
  2347 => x"c002bfc4",
  2348 => x"c14887c9",
  2349 => x"c8f4c288",
  2350 => x"c487d358",
  2351 => x"e0c14866",
  2352 => x"6e7e7080",
  2353 => x"c5c002bf",
  2354 => x"49ff4b87",
  2355 => x"a6c80f73",
  2356 => x"7478c148",
  2357 => x"0599c449",
  2358 => x"c387cec0",
  2359 => x"fae249f2",
  2360 => x"c2497087",
  2361 => x"f0c00299",
  2362 => x"c4f4c287",
  2363 => x"c7487ebf",
  2364 => x"c003a8b7",
  2365 => x"486e87cb",
  2366 => x"f4c280c1",
  2367 => x"d3c058c8",
  2368 => x"4866c487",
  2369 => x"7080e0c1",
  2370 => x"02bf6e7e",
  2371 => x"4b87c5c0",
  2372 => x"0f7349fe",
  2373 => x"c148a6c8",
  2374 => x"49fdc378",
  2375 => x"7087fce1",
  2376 => x"0299c249",
  2377 => x"c287e9c0",
  2378 => x"02bfc4f4",
  2379 => x"c287c9c0",
  2380 => x"c048c4f4",
  2381 => x"87d3c078",
  2382 => x"c14866c4",
  2383 => x"7e7080e0",
  2384 => x"c002bf6e",
  2385 => x"fd4b87c5",
  2386 => x"c80f7349",
  2387 => x"78c148a6",
  2388 => x"e149fac3",
  2389 => x"497087c5",
  2390 => x"c00299c2",
  2391 => x"f4c287ea",
  2392 => x"c748bfc4",
  2393 => x"c003a8b7",
  2394 => x"f4c287c9",
  2395 => x"78c748c4",
  2396 => x"c487d0c0",
  2397 => x"e0c14a66",
  2398 => x"c0026a82",
  2399 => x"fc4b87c5",
  2400 => x"c80f7349",
  2401 => x"78c148a6",
  2402 => x"f3c24dc0",
  2403 => x"50c048fc",
  2404 => x"c249eecb",
  2405 => x"4b7087f2",
  2406 => x"97fcf3c2",
  2407 => x"ddc105bf",
  2408 => x"c3497487",
  2409 => x"c00599f0",
  2410 => x"dac187cd",
  2411 => x"eadfff49",
  2412 => x"02987087",
  2413 => x"c187c7c1",
  2414 => x"4cbfe84d",
  2415 => x"99ffc349",
  2416 => x"712cb7c8",
  2417 => x"c4d9c2b4",
  2418 => x"dbff49bf",
  2419 => x"497387cb",
  2420 => x"7087c1c2",
  2421 => x"c6c00298",
  2422 => x"fcf3c287",
  2423 => x"c250c148",
  2424 => x"bf97fcf3",
  2425 => x"87d6c005",
  2426 => x"f0c34974",
  2427 => x"c6ff0599",
  2428 => x"49dac187",
  2429 => x"87e3deff",
  2430 => x"fe059870",
  2431 => x"9d7587f9",
  2432 => x"87e0c002",
  2433 => x"c248a6cc",
  2434 => x"78bfc4f4",
  2435 => x"cc4966cc",
  2436 => x"4866c491",
  2437 => x"7e708071",
  2438 => x"c002bf6e",
  2439 => x"cc4b87c6",
  2440 => x"0f734966",
  2441 => x"c00266c8",
  2442 => x"f4c287c8",
  2443 => x"f249bfc4",
  2444 => x"8ef087ce",
  2445 => x"4c264d26",
  2446 => x"4f264b26",
  2447 => x"00000000",
  2448 => x"00000000",
  2449 => x"00000000",
  2450 => x"ff4a711e",
  2451 => x"7249bfc8",
  2452 => x"4f2648a1",
  2453 => x"bfc8ff1e",
  2454 => x"c0c0fe89",
  2455 => x"a9c0c0c0",
  2456 => x"c087c401",
  2457 => x"c187c24a",
  2458 => x"2648724a",
  2459 => x"5b5e0e4f",
  2460 => x"710e5d5c",
  2461 => x"4cd4ff4b",
  2462 => x"c04866d0",
  2463 => x"ff49d678",
  2464 => x"c387d5de",
  2465 => x"496c7cff",
  2466 => x"7199ffc3",
  2467 => x"f0c3494d",
  2468 => x"a9e0c199",
  2469 => x"c387cb05",
  2470 => x"486c7cff",
  2471 => x"66d098c3",
  2472 => x"ffc37808",
  2473 => x"494a6c7c",
  2474 => x"ffc331c8",
  2475 => x"714a6c7c",
  2476 => x"c84972b2",
  2477 => x"7cffc331",
  2478 => x"b2714a6c",
  2479 => x"31c84972",
  2480 => x"6c7cffc3",
  2481 => x"ffb2714a",
  2482 => x"e0c048d0",
  2483 => x"029b7378",
  2484 => x"7b7287c2",
  2485 => x"4d264875",
  2486 => x"4b264c26",
  2487 => x"261e4f26",
  2488 => x"5b5e0e4f",
  2489 => x"86f80e5c",
  2490 => x"a6c81e76",
  2491 => x"87fdfd49",
  2492 => x"4b7086c4",
  2493 => x"a8c2486e",
  2494 => x"87f0c203",
  2495 => x"f0c34a73",
  2496 => x"aad0c19a",
  2497 => x"c187c702",
  2498 => x"c205aae0",
  2499 => x"497387de",
  2500 => x"c30299c8",
  2501 => x"87c6ff87",
  2502 => x"9cc34c73",
  2503 => x"c105acc2",
  2504 => x"66c487c2",
  2505 => x"7131c949",
  2506 => x"4a66c41e",
  2507 => x"f4c292d4",
  2508 => x"817249c8",
  2509 => x"87dccefe",
  2510 => x"dbff49d8",
  2511 => x"c0c887da",
  2512 => x"e0e2c21e",
  2513 => x"cee8fd49",
  2514 => x"48d0ff87",
  2515 => x"c278e0c0",
  2516 => x"cc1ee0e2",
  2517 => x"92d44a66",
  2518 => x"49c8f4c2",
  2519 => x"ccfe8172",
  2520 => x"86cc87e3",
  2521 => x"c105acc1",
  2522 => x"66c487c2",
  2523 => x"7131c949",
  2524 => x"4a66c41e",
  2525 => x"f4c292d4",
  2526 => x"817249c8",
  2527 => x"87d4cdfe",
  2528 => x"1ee0e2c2",
  2529 => x"d44a66c8",
  2530 => x"c8f4c292",
  2531 => x"fe817249",
  2532 => x"d787e3ca",
  2533 => x"ffd9ff49",
  2534 => x"1ec0c887",
  2535 => x"49e0e2c2",
  2536 => x"87d0e6fd",
  2537 => x"d0ff86cc",
  2538 => x"78e0c048",
  2539 => x"4c268ef8",
  2540 => x"4f264b26",
  2541 => x"5c5b5e0e",
  2542 => x"86fc0e5d",
  2543 => x"d4ff4d71",
  2544 => x"7e66d44c",
  2545 => x"a8b7c348",
  2546 => x"87e2c101",
  2547 => x"66c41e75",
  2548 => x"c293d44b",
  2549 => x"7383c8f4",
  2550 => x"d8c4fe49",
  2551 => x"49a3c887",
  2552 => x"d0ff4969",
  2553 => x"78e1c848",
  2554 => x"48717cdd",
  2555 => x"7098ffc3",
  2556 => x"c84a717c",
  2557 => x"48722ab7",
  2558 => x"7098ffc3",
  2559 => x"d04a717c",
  2560 => x"48722ab7",
  2561 => x"7098ffc3",
  2562 => x"d848717c",
  2563 => x"7c7028b7",
  2564 => x"7c7c7cc0",
  2565 => x"7c7c7c7c",
  2566 => x"7c7c7c7c",
  2567 => x"48d0ff7c",
  2568 => x"c478e0c0",
  2569 => x"49dc1e66",
  2570 => x"87d1d8ff",
  2571 => x"8efc86c8",
  2572 => x"4c264d26",
  2573 => x"4f264b26",
  2574 => x"c21ec01e",
  2575 => x"49bfd4e1",
  2576 => x"c287f1fd",
  2577 => x"49bfd8e1",
  2578 => x"87fadcfe",
  2579 => x"8efc48c0",
  2580 => x"00004f26",
  2581 => x"0000285c",
  2582 => x"00002868",
  2583 => x"20434242",
  2584 => x"20202020",
  2585 => x"00444856",
  2586 => x"20434242",
  2587 => x"20202020",
  2588 => x"004d4f52",
  2589 => x"00001baf",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
