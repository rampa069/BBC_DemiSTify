library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d0efc287",
    12 => x"86c0c84e",
    13 => x"49d0efc2",
    14 => x"48e8dcc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087f2df",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d40299",
    50 => x"d4ff4812",
    51 => x"66c47808",
    52 => x"88c14849",
    53 => x"7158a6c8",
    54 => x"87ec0599",
    55 => x"711e4f26",
    56 => x"4966c44a",
    57 => x"c888c148",
    58 => x"997158a6",
    59 => x"ff87d602",
    60 => x"ffc348d4",
    61 => x"c4526878",
    62 => x"c1484966",
    63 => x"58a6c888",
    64 => x"ea059971",
    65 => x"1e4f2687",
    66 => x"d4ff1e73",
    67 => x"7bffc34b",
    68 => x"ffc34a6b",
    69 => x"c8496b7b",
    70 => x"c3b17232",
    71 => x"4a6b7bff",
    72 => x"b27131c8",
    73 => x"6b7bffc3",
    74 => x"7232c849",
    75 => x"c44871b1",
    76 => x"264d2687",
    77 => x"264b264c",
    78 => x"5b5e0e4f",
    79 => x"710e5d5c",
    80 => x"4cd4ff4a",
    81 => x"ffc34872",
    82 => x"c27c7098",
    83 => x"05bfe8dc",
    84 => x"66d087c8",
    85 => x"d430c948",
    86 => x"66d058a6",
    87 => x"7129d849",
    88 => x"98ffc348",
    89 => x"66d07c70",
    90 => x"7129d049",
    91 => x"98ffc348",
    92 => x"66d07c70",
    93 => x"7129c849",
    94 => x"98ffc348",
    95 => x"66d07c70",
    96 => x"98ffc348",
    97 => x"49727c70",
    98 => x"487129d0",
    99 => x"7098ffc3",
   100 => x"c94b6c7c",
   101 => x"c34dfff0",
   102 => x"d005abff",
   103 => x"7cffc387",
   104 => x"8dc14b6c",
   105 => x"c387c602",
   106 => x"f002abff",
   107 => x"fd487387",
   108 => x"c01e87ff",
   109 => x"48d4ff49",
   110 => x"c178ffc3",
   111 => x"b7c8c381",
   112 => x"87f104a9",
   113 => x"731e4f26",
   114 => x"c487e71e",
   115 => x"c04bdff8",
   116 => x"f0ffc01e",
   117 => x"fd49f7c1",
   118 => x"86c487df",
   119 => x"c005a8c1",
   120 => x"d4ff87ea",
   121 => x"78ffc348",
   122 => x"c0c0c0c1",
   123 => x"c01ec0c0",
   124 => x"e9c1f0e1",
   125 => x"87c1fd49",
   126 => x"987086c4",
   127 => x"ff87ca05",
   128 => x"ffc348d4",
   129 => x"cb48c178",
   130 => x"87e6fe87",
   131 => x"fe058bc1",
   132 => x"48c087fd",
   133 => x"1e87defc",
   134 => x"d4ff1e73",
   135 => x"78ffc348",
   136 => x"1ec04bd3",
   137 => x"c1f0ffc0",
   138 => x"ccfc49c1",
   139 => x"7086c487",
   140 => x"87ca0598",
   141 => x"c348d4ff",
   142 => x"48c178ff",
   143 => x"f1fd87cb",
   144 => x"058bc187",
   145 => x"c087dbff",
   146 => x"87e9fb48",
   147 => x"5c5b5e0e",
   148 => x"4cd4ff0e",
   149 => x"c687dbfd",
   150 => x"e1c01eea",
   151 => x"49c8c1f0",
   152 => x"c487d6fb",
   153 => x"02a8c186",
   154 => x"eafe87c8",
   155 => x"c148c087",
   156 => x"d2fa87e2",
   157 => x"cf497087",
   158 => x"c699ffff",
   159 => x"c802a9ea",
   160 => x"87d3fe87",
   161 => x"cbc148c0",
   162 => x"7cffc387",
   163 => x"fc4bf1c0",
   164 => x"987087f4",
   165 => x"87ebc002",
   166 => x"ffc01ec0",
   167 => x"49fac1f0",
   168 => x"c487d6fa",
   169 => x"05987086",
   170 => x"ffc387d9",
   171 => x"c3496c7c",
   172 => x"7c7c7cff",
   173 => x"99c0c17c",
   174 => x"c187c402",
   175 => x"c087d548",
   176 => x"c287d148",
   177 => x"87c405ab",
   178 => x"87c848c0",
   179 => x"fe058bc1",
   180 => x"48c087fd",
   181 => x"1e87dcf9",
   182 => x"dcc21e73",
   183 => x"78c148e8",
   184 => x"d0ff4bc7",
   185 => x"fb78c248",
   186 => x"d0ff87c8",
   187 => x"c078c348",
   188 => x"d0e5c01e",
   189 => x"f849c0c1",
   190 => x"86c487ff",
   191 => x"c105a8c1",
   192 => x"abc24b87",
   193 => x"c087c505",
   194 => x"87f9c048",
   195 => x"ff058bc1",
   196 => x"f7fc87d0",
   197 => x"ecdcc287",
   198 => x"05987058",
   199 => x"1ec187cd",
   200 => x"c1f0ffc0",
   201 => x"d0f849d0",
   202 => x"ff86c487",
   203 => x"ffc348d4",
   204 => x"87ddc478",
   205 => x"58f0dcc2",
   206 => x"c248d0ff",
   207 => x"48d4ff78",
   208 => x"c178ffc3",
   209 => x"87edf748",
   210 => x"5c5b5e0e",
   211 => x"4a710e5d",
   212 => x"ff4dffc3",
   213 => x"7c754cd4",
   214 => x"c448d0ff",
   215 => x"7c7578c3",
   216 => x"ffc01e72",
   217 => x"49d8c1f0",
   218 => x"c487cef7",
   219 => x"02987086",
   220 => x"48c187c5",
   221 => x"7587eec0",
   222 => x"7cfec37c",
   223 => x"d41ec0c8",
   224 => x"f2f44966",
   225 => x"7586c487",
   226 => x"757c757c",
   227 => x"e0dad87c",
   228 => x"6c7c754b",
   229 => x"c187c505",
   230 => x"87f5058b",
   231 => x"d0ff7c75",
   232 => x"c078c248",
   233 => x"87c9f648",
   234 => x"5c5b5e0e",
   235 => x"4b710e5d",
   236 => x"eec54cc0",
   237 => x"ff4adfcd",
   238 => x"ffc348d4",
   239 => x"c3486878",
   240 => x"c005a8fe",
   241 => x"d4ff87fe",
   242 => x"029b734d",
   243 => x"66d087cc",
   244 => x"f449731e",
   245 => x"86c487c8",
   246 => x"d0ff87d6",
   247 => x"78d1c448",
   248 => x"d07dffc3",
   249 => x"88c14866",
   250 => x"7058a6d4",
   251 => x"87f00598",
   252 => x"c348d4ff",
   253 => x"737878ff",
   254 => x"87c5059b",
   255 => x"d048d0ff",
   256 => x"4c4ac178",
   257 => x"fe058ac1",
   258 => x"487487ed",
   259 => x"1e87e2f4",
   260 => x"4a711e73",
   261 => x"d4ff4bc0",
   262 => x"78ffc348",
   263 => x"c448d0ff",
   264 => x"d4ff78c3",
   265 => x"78ffc348",
   266 => x"ffc01e72",
   267 => x"49d1c1f0",
   268 => x"c487c6f4",
   269 => x"05987086",
   270 => x"c0c887d2",
   271 => x"4966cc1e",
   272 => x"c487e5fd",
   273 => x"ff4b7086",
   274 => x"78c248d0",
   275 => x"e4f34873",
   276 => x"5b5e0e87",
   277 => x"c00e5d5c",
   278 => x"f0ffc01e",
   279 => x"f349c9c1",
   280 => x"1ed287d7",
   281 => x"49f0dcc2",
   282 => x"c887fdfc",
   283 => x"c14cc086",
   284 => x"acb7d284",
   285 => x"c287f804",
   286 => x"bf97f0dc",
   287 => x"99c0c349",
   288 => x"05a9c0c1",
   289 => x"c287e7c0",
   290 => x"bf97f7dc",
   291 => x"c231d049",
   292 => x"bf97f8dc",
   293 => x"7232c84a",
   294 => x"f9dcc2b1",
   295 => x"b14abf97",
   296 => x"ffcf4c71",
   297 => x"c19cffff",
   298 => x"c134ca84",
   299 => x"dcc287e7",
   300 => x"49bf97f9",
   301 => x"99c631c1",
   302 => x"97fadcc2",
   303 => x"b7c74abf",
   304 => x"c2b1722a",
   305 => x"bf97f5dc",
   306 => x"9dcf4d4a",
   307 => x"97f6dcc2",
   308 => x"9ac34abf",
   309 => x"dcc232ca",
   310 => x"4bbf97f7",
   311 => x"b27333c2",
   312 => x"97f8dcc2",
   313 => x"c0c34bbf",
   314 => x"2bb7c69b",
   315 => x"81c2b273",
   316 => x"307148c1",
   317 => x"48c14970",
   318 => x"4d703075",
   319 => x"84c14c72",
   320 => x"c0c89471",
   321 => x"cc06adb7",
   322 => x"b734c187",
   323 => x"b7c0c82d",
   324 => x"f4ff01ad",
   325 => x"f0487487",
   326 => x"5e0e87d7",
   327 => x"0e5d5c5b",
   328 => x"e5c286f8",
   329 => x"78c048d6",
   330 => x"1eceddc2",
   331 => x"defb49c0",
   332 => x"7086c487",
   333 => x"87c50598",
   334 => x"c0c948c0",
   335 => x"c14dc087",
   336 => x"ddf2c07e",
   337 => x"dec249bf",
   338 => x"c8714ac4",
   339 => x"87d9ec4b",
   340 => x"c2059870",
   341 => x"c07ec087",
   342 => x"49bfd9f2",
   343 => x"4ae0dec2",
   344 => x"ec4bc871",
   345 => x"987087c3",
   346 => x"c087c205",
   347 => x"c0026e7e",
   348 => x"e4c287fd",
   349 => x"c24dbfd4",
   350 => x"bf9fcce5",
   351 => x"d6c5487e",
   352 => x"c705a8ea",
   353 => x"d4e4c287",
   354 => x"87ce4dbf",
   355 => x"e9ca486e",
   356 => x"c502a8d5",
   357 => x"c748c087",
   358 => x"ddc287e3",
   359 => x"49751ece",
   360 => x"c487ecf9",
   361 => x"05987086",
   362 => x"48c087c5",
   363 => x"c087cec7",
   364 => x"49bfd9f2",
   365 => x"4ae0dec2",
   366 => x"ea4bc871",
   367 => x"987087eb",
   368 => x"c287c805",
   369 => x"c148d6e5",
   370 => x"c087da78",
   371 => x"49bfddf2",
   372 => x"4ac4dec2",
   373 => x"ea4bc871",
   374 => x"987087cf",
   375 => x"87c5c002",
   376 => x"d8c648c0",
   377 => x"cce5c287",
   378 => x"c149bf97",
   379 => x"c005a9d5",
   380 => x"e5c287cd",
   381 => x"49bf97cd",
   382 => x"02a9eac2",
   383 => x"c087c5c0",
   384 => x"87f9c548",
   385 => x"97ceddc2",
   386 => x"c3487ebf",
   387 => x"c002a8e9",
   388 => x"486e87ce",
   389 => x"02a8ebc3",
   390 => x"c087c5c0",
   391 => x"87ddc548",
   392 => x"97d9ddc2",
   393 => x"059949bf",
   394 => x"c287ccc0",
   395 => x"bf97dadd",
   396 => x"02a9c249",
   397 => x"c087c5c0",
   398 => x"87c1c548",
   399 => x"97dbddc2",
   400 => x"e5c248bf",
   401 => x"4c7058d2",
   402 => x"c288c148",
   403 => x"c258d6e5",
   404 => x"bf97dcdd",
   405 => x"c2817549",
   406 => x"bf97dddd",
   407 => x"7232c84a",
   408 => x"e9c27ea1",
   409 => x"786e48e3",
   410 => x"97deddc2",
   411 => x"a6c848bf",
   412 => x"d6e5c258",
   413 => x"cfc202bf",
   414 => x"d9f2c087",
   415 => x"dec249bf",
   416 => x"c8714ae0",
   417 => x"87e1e74b",
   418 => x"c0029870",
   419 => x"48c087c5",
   420 => x"c287eac3",
   421 => x"4cbfcee5",
   422 => x"5cf7e9c2",
   423 => x"97f3ddc2",
   424 => x"31c849bf",
   425 => x"97f2ddc2",
   426 => x"49a14abf",
   427 => x"97f4ddc2",
   428 => x"32d04abf",
   429 => x"c249a172",
   430 => x"bf97f5dd",
   431 => x"7232d84a",
   432 => x"66c449a1",
   433 => x"e3e9c291",
   434 => x"e9c281bf",
   435 => x"ddc259eb",
   436 => x"4abf97fb",
   437 => x"ddc232c8",
   438 => x"4bbf97fa",
   439 => x"ddc24aa2",
   440 => x"4bbf97fc",
   441 => x"a27333d0",
   442 => x"fdddc24a",
   443 => x"cf4bbf97",
   444 => x"7333d89b",
   445 => x"e9c24aa2",
   446 => x"8ac25aef",
   447 => x"e9c29274",
   448 => x"a17248ef",
   449 => x"87c1c178",
   450 => x"97e0ddc2",
   451 => x"31c849bf",
   452 => x"97dfddc2",
   453 => x"49a14abf",
   454 => x"ffc731c5",
   455 => x"c229c981",
   456 => x"c259f7e9",
   457 => x"bf97e5dd",
   458 => x"c232c84a",
   459 => x"bf97e4dd",
   460 => x"c44aa24b",
   461 => x"826e9266",
   462 => x"5af3e9c2",
   463 => x"48ebe9c2",
   464 => x"e9c278c0",
   465 => x"a17248e7",
   466 => x"f7e9c278",
   467 => x"ebe9c248",
   468 => x"e9c278bf",
   469 => x"e9c248fb",
   470 => x"c278bfef",
   471 => x"02bfd6e5",
   472 => x"7487c9c0",
   473 => x"7030c448",
   474 => x"87c9c07e",
   475 => x"bff3e9c2",
   476 => x"7030c448",
   477 => x"dae5c27e",
   478 => x"c1786e48",
   479 => x"268ef848",
   480 => x"264c264d",
   481 => x"0e4f264b",
   482 => x"5d5c5b5e",
   483 => x"c24a710e",
   484 => x"02bfd6e5",
   485 => x"4b7287cb",
   486 => x"4d722bc7",
   487 => x"c99dffc1",
   488 => x"c84b7287",
   489 => x"c34d722b",
   490 => x"e9c29dff",
   491 => x"c083bfe3",
   492 => x"abbfd5f2",
   493 => x"c087d902",
   494 => x"c25bd9f2",
   495 => x"731ecedd",
   496 => x"87cbf149",
   497 => x"987086c4",
   498 => x"c087c505",
   499 => x"87e6c048",
   500 => x"bfd6e5c2",
   501 => x"7587d202",
   502 => x"c291c449",
   503 => x"6981cedd",
   504 => x"ffffcf4c",
   505 => x"cb9cffff",
   506 => x"c2497587",
   507 => x"ceddc291",
   508 => x"4c699f81",
   509 => x"c6fe4874",
   510 => x"5b5e0e87",
   511 => x"f80e5d5c",
   512 => x"9c4c7186",
   513 => x"c087c505",
   514 => x"87c0c348",
   515 => x"487ea4c8",
   516 => x"66d878c0",
   517 => x"d887c702",
   518 => x"05bf9766",
   519 => x"48c087c5",
   520 => x"c087e9c2",
   521 => x"4949c11e",
   522 => x"c487d3ca",
   523 => x"9d4d7086",
   524 => x"87c2c102",
   525 => x"4adee5c2",
   526 => x"e04966d8",
   527 => x"987087d0",
   528 => x"87f2c002",
   529 => x"66d84a75",
   530 => x"e04bcb49",
   531 => x"987087f5",
   532 => x"87e2c002",
   533 => x"9d751ec0",
   534 => x"c887c702",
   535 => x"78c048a6",
   536 => x"a6c887c5",
   537 => x"c878c148",
   538 => x"d1c94966",
   539 => x"7086c487",
   540 => x"fe059d4d",
   541 => x"9d7587fe",
   542 => x"87cec102",
   543 => x"6e49a5dc",
   544 => x"da786948",
   545 => x"a6c449a5",
   546 => x"78a4c448",
   547 => x"c448699f",
   548 => x"c2780866",
   549 => x"02bfd6e5",
   550 => x"a5d487d2",
   551 => x"49699f49",
   552 => x"99ffffc0",
   553 => x"30d04871",
   554 => x"87c27e70",
   555 => x"486e7ec0",
   556 => x"80bf66c4",
   557 => x"780866c4",
   558 => x"a4cc7cc0",
   559 => x"bf66c449",
   560 => x"49a4d079",
   561 => x"48c179c0",
   562 => x"48c087c2",
   563 => x"eefa8ef8",
   564 => x"5b5e0e87",
   565 => x"4c710e5c",
   566 => x"cbc1029c",
   567 => x"49a4c887",
   568 => x"c3c10269",
   569 => x"cc496c87",
   570 => x"80714866",
   571 => x"7058a6d0",
   572 => x"d2e5c2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e5c002",
   576 => x"6b4ba4c4",
   577 => x"87fff949",
   578 => x"e5c27b70",
   579 => x"6c49bfce",
   580 => x"cc7c7181",
   581 => x"e5c2b966",
   582 => x"ff4abfd2",
   583 => x"719972ba",
   584 => x"dbff0599",
   585 => x"7c66cc87",
   586 => x"1e87d6f9",
   587 => x"4b711e73",
   588 => x"87c7029b",
   589 => x"6949a3c8",
   590 => x"c087c505",
   591 => x"87f6c048",
   592 => x"bfe7e9c2",
   593 => x"4aa3c449",
   594 => x"8ac24a6a",
   595 => x"bfcee5c2",
   596 => x"49a17292",
   597 => x"bfd2e5c2",
   598 => x"729a6b4a",
   599 => x"f2c049a1",
   600 => x"66c859d9",
   601 => x"e6ea711e",
   602 => x"7086c487",
   603 => x"87c40598",
   604 => x"87c248c0",
   605 => x"caf848c1",
   606 => x"1e731e87",
   607 => x"029b4b71",
   608 => x"a3c887c7",
   609 => x"c5056949",
   610 => x"c048c087",
   611 => x"e9c287f6",
   612 => x"c449bfe7",
   613 => x"4a6a4aa3",
   614 => x"e5c28ac2",
   615 => x"7292bfce",
   616 => x"e5c249a1",
   617 => x"6b4abfd2",
   618 => x"49a1729a",
   619 => x"59d9f2c0",
   620 => x"711e66c8",
   621 => x"c487d1e6",
   622 => x"05987086",
   623 => x"48c087c4",
   624 => x"48c187c2",
   625 => x"0e87fcf6",
   626 => x"5d5c5b5e",
   627 => x"4b711e0e",
   628 => x"734d66d4",
   629 => x"ccc1029b",
   630 => x"49a3c887",
   631 => x"c4c10269",
   632 => x"4ca3d087",
   633 => x"bfd2e5c2",
   634 => x"6cb9ff49",
   635 => x"d47e994a",
   636 => x"cd06a966",
   637 => x"7c7bc087",
   638 => x"c44aa3cc",
   639 => x"796a49a3",
   640 => x"497287ca",
   641 => x"d499c0f8",
   642 => x"8d714d66",
   643 => x"29c94975",
   644 => x"49731e71",
   645 => x"c287fafa",
   646 => x"731ecedd",
   647 => x"87cbfc49",
   648 => x"66d486c8",
   649 => x"d6f5267c",
   650 => x"1e731e87",
   651 => x"029b4b71",
   652 => x"c287e4c0",
   653 => x"735bfbe9",
   654 => x"c28ac24a",
   655 => x"49bfcee5",
   656 => x"e7e9c292",
   657 => x"807248bf",
   658 => x"58ffe9c2",
   659 => x"30c44871",
   660 => x"58dee5c2",
   661 => x"c287edc0",
   662 => x"c248f7e9",
   663 => x"78bfebe9",
   664 => x"48fbe9c2",
   665 => x"bfefe9c2",
   666 => x"d6e5c278",
   667 => x"87c902bf",
   668 => x"bfcee5c2",
   669 => x"c731c449",
   670 => x"f3e9c287",
   671 => x"31c449bf",
   672 => x"59dee5c2",
   673 => x"0e87fcf3",
   674 => x"0e5c5b5e",
   675 => x"4bc04a71",
   676 => x"c0029a72",
   677 => x"a2da87e0",
   678 => x"4b699f49",
   679 => x"bfd6e5c2",
   680 => x"d487cf02",
   681 => x"699f49a2",
   682 => x"ffc04c49",
   683 => x"34d09cff",
   684 => x"4cc087c2",
   685 => x"4973b374",
   686 => x"f387eefd",
   687 => x"5e0e87c3",
   688 => x"0e5d5c5b",
   689 => x"4a7186f4",
   690 => x"9a727ec0",
   691 => x"c287d802",
   692 => x"c048cadd",
   693 => x"c2ddc278",
   694 => x"fbe9c248",
   695 => x"ddc278bf",
   696 => x"e9c248c6",
   697 => x"c278bff7",
   698 => x"c048ebe5",
   699 => x"dae5c250",
   700 => x"ddc249bf",
   701 => x"714abfca",
   702 => x"c9c403aa",
   703 => x"cf497287",
   704 => x"e9c00599",
   705 => x"d5f2c087",
   706 => x"c2ddc248",
   707 => x"ddc278bf",
   708 => x"ddc21ece",
   709 => x"c249bfc2",
   710 => x"c148c2dd",
   711 => x"e37178a1",
   712 => x"86c487ed",
   713 => x"48d1f2c0",
   714 => x"78ceddc2",
   715 => x"f2c087cc",
   716 => x"c048bfd1",
   717 => x"f2c080e0",
   718 => x"ddc258d5",
   719 => x"c148bfca",
   720 => x"ceddc280",
   721 => x"0c912758",
   722 => x"97bf0000",
   723 => x"029d4dbf",
   724 => x"c387e3c2",
   725 => x"c202ade5",
   726 => x"f2c087dc",
   727 => x"cb4bbfd1",
   728 => x"4c1149a3",
   729 => x"c105accf",
   730 => x"497587d2",
   731 => x"89c199df",
   732 => x"e5c291cd",
   733 => x"a3c181de",
   734 => x"c351124a",
   735 => x"51124aa3",
   736 => x"124aa3c5",
   737 => x"4aa3c751",
   738 => x"a3c95112",
   739 => x"ce51124a",
   740 => x"51124aa3",
   741 => x"124aa3d0",
   742 => x"4aa3d251",
   743 => x"a3d45112",
   744 => x"d651124a",
   745 => x"51124aa3",
   746 => x"124aa3d8",
   747 => x"4aa3dc51",
   748 => x"a3de5112",
   749 => x"c151124a",
   750 => x"87fac07e",
   751 => x"99c84974",
   752 => x"87ebc005",
   753 => x"99d04974",
   754 => x"dc87d105",
   755 => x"cbc00266",
   756 => x"dc497387",
   757 => x"98700f66",
   758 => x"87d3c002",
   759 => x"c6c0056e",
   760 => x"dee5c287",
   761 => x"c050c048",
   762 => x"48bfd1f2",
   763 => x"c287ddc2",
   764 => x"c048ebe5",
   765 => x"e5c27e50",
   766 => x"c249bfda",
   767 => x"4abfcadd",
   768 => x"fb04aa71",
   769 => x"e9c287f7",
   770 => x"c005bffb",
   771 => x"e5c287c8",
   772 => x"c102bfd6",
   773 => x"ddc287f4",
   774 => x"ed49bfc6",
   775 => x"ddc287e9",
   776 => x"a6c458ca",
   777 => x"c6ddc248",
   778 => x"e5c278bf",
   779 => x"c002bfd6",
   780 => x"66c487d8",
   781 => x"ffffcf49",
   782 => x"a999f8ff",
   783 => x"87c5c002",
   784 => x"e1c04cc0",
   785 => x"c04cc187",
   786 => x"66c487dc",
   787 => x"f8ffcf49",
   788 => x"c002a999",
   789 => x"a6c887c8",
   790 => x"c078c048",
   791 => x"a6c887c5",
   792 => x"c878c148",
   793 => x"9c744c66",
   794 => x"87dec005",
   795 => x"c24966c4",
   796 => x"cee5c289",
   797 => x"e9c291bf",
   798 => x"7148bfe7",
   799 => x"c6ddc280",
   800 => x"caddc258",
   801 => x"f978c048",
   802 => x"48c087e3",
   803 => x"eeeb8ef4",
   804 => x"00000087",
   805 => x"ffffff00",
   806 => x"000ca1ff",
   807 => x"000caa00",
   808 => x"54414600",
   809 => x"20203233",
   810 => x"41460020",
   811 => x"20363154",
   812 => x"1e002020",
   813 => x"c348d4ff",
   814 => x"486878ff",
   815 => x"ff1e4f26",
   816 => x"ffc348d4",
   817 => x"48d0ff78",
   818 => x"ff78e1c0",
   819 => x"78d448d4",
   820 => x"48ffe9c2",
   821 => x"50bfd4ff",
   822 => x"ff1e4f26",
   823 => x"e0c048d0",
   824 => x"1e4f2678",
   825 => x"7087ccff",
   826 => x"c6029949",
   827 => x"a9fbc087",
   828 => x"7187f105",
   829 => x"0e4f2648",
   830 => x"0e5c5b5e",
   831 => x"4cc04b71",
   832 => x"7087f0fe",
   833 => x"c0029949",
   834 => x"ecc087f9",
   835 => x"f2c002a9",
   836 => x"a9fbc087",
   837 => x"87ebc002",
   838 => x"acb766cc",
   839 => x"d087c703",
   840 => x"87c20266",
   841 => x"99715371",
   842 => x"c187c202",
   843 => x"87c3fe84",
   844 => x"02994970",
   845 => x"ecc087cd",
   846 => x"87c702a9",
   847 => x"05a9fbc0",
   848 => x"d087d5ff",
   849 => x"87c30266",
   850 => x"c07b97c0",
   851 => x"c405a9ec",
   852 => x"c54a7487",
   853 => x"c04a7487",
   854 => x"48728a0a",
   855 => x"4d2687c2",
   856 => x"4b264c26",
   857 => x"fd1e4f26",
   858 => x"497087c9",
   859 => x"aaf0c04a",
   860 => x"c087c904",
   861 => x"c301aaf9",
   862 => x"8af0c087",
   863 => x"04aac1c1",
   864 => x"dac187c9",
   865 => x"87c301aa",
   866 => x"728af7c0",
   867 => x"0e4f2648",
   868 => x"5d5c5b5e",
   869 => x"7186f80e",
   870 => x"fc4dc04c",
   871 => x"4bc087e0",
   872 => x"97eef8c0",
   873 => x"a9c049bf",
   874 => x"fc87cf04",
   875 => x"83c187f5",
   876 => x"97eef8c0",
   877 => x"06ab49bf",
   878 => x"f8c087f1",
   879 => x"02bf97ee",
   880 => x"eefb87cf",
   881 => x"99497087",
   882 => x"c087c602",
   883 => x"f105a9ec",
   884 => x"fb4bc087",
   885 => x"7e7087dd",
   886 => x"c887d8fb",
   887 => x"d2fb58a6",
   888 => x"c14a7087",
   889 => x"49a4c883",
   890 => x"6e496997",
   891 => x"87da05a9",
   892 => x"9749a4c9",
   893 => x"66c44969",
   894 => x"87ce05a9",
   895 => x"9749a4ca",
   896 => x"05aa4969",
   897 => x"4dc187c4",
   898 => x"486e87d4",
   899 => x"02a8ecc0",
   900 => x"486e87c8",
   901 => x"05a8fbc0",
   902 => x"4bc087c4",
   903 => x"9d754dc1",
   904 => x"87effe02",
   905 => x"7387f3fa",
   906 => x"fc8ef848",
   907 => x"0e0087f0",
   908 => x"5d5c5b5e",
   909 => x"7186f80e",
   910 => x"4bd4ff7e",
   911 => x"eac21e6e",
   912 => x"f4e649c4",
   913 => x"7086c487",
   914 => x"eac40298",
   915 => x"c2e3c187",
   916 => x"496e4dbf",
   917 => x"c887f8fc",
   918 => x"987058a6",
   919 => x"c487c505",
   920 => x"78c148a6",
   921 => x"c548d0ff",
   922 => x"7bd5c178",
   923 => x"c14966c4",
   924 => x"c131c689",
   925 => x"bf97c0e3",
   926 => x"b071484a",
   927 => x"d0ff7b70",
   928 => x"c278c448",
   929 => x"bf97ffe9",
   930 => x"0299d049",
   931 => x"78c587d7",
   932 => x"c07bd6c1",
   933 => x"7bffc34a",
   934 => x"e0c082c1",
   935 => x"87f504aa",
   936 => x"c448d0ff",
   937 => x"7bffc378",
   938 => x"c548d0ff",
   939 => x"7bd3c178",
   940 => x"78c47bc1",
   941 => x"06adb7c0",
   942 => x"c287ebc2",
   943 => x"4cbfccea",
   944 => x"c2029c8d",
   945 => x"ddc287c2",
   946 => x"a6c47ece",
   947 => x"78c0c848",
   948 => x"acb7c08c",
   949 => x"c887c603",
   950 => x"c078a4c0",
   951 => x"ffe9c24c",
   952 => x"d049bf97",
   953 => x"87d00299",
   954 => x"eac21ec0",
   955 => x"fae849c4",
   956 => x"7086c487",
   957 => x"87f5c04a",
   958 => x"1eceddc2",
   959 => x"49c4eac2",
   960 => x"c487e8e8",
   961 => x"ff4a7086",
   962 => x"c5c848d0",
   963 => x"7bd4c178",
   964 => x"7bbf976e",
   965 => x"80c1486e",
   966 => x"66c47e70",
   967 => x"c888c148",
   968 => x"987058a6",
   969 => x"87e8ff05",
   970 => x"c448d0ff",
   971 => x"059a7278",
   972 => x"48c087c5",
   973 => x"c187c2c1",
   974 => x"c4eac21e",
   975 => x"87d1e649",
   976 => x"9c7486c4",
   977 => x"87fefd05",
   978 => x"06adb7c0",
   979 => x"eac287d1",
   980 => x"78c048c4",
   981 => x"78c080d0",
   982 => x"eac280f4",
   983 => x"c078bfd0",
   984 => x"fd01adb7",
   985 => x"d0ff87d5",
   986 => x"c178c548",
   987 => x"7bc07bd3",
   988 => x"48c178c4",
   989 => x"c087c2c0",
   990 => x"268ef848",
   991 => x"264c264d",
   992 => x"0e4f264b",
   993 => x"5d5c5b5e",
   994 => x"4b711e0e",
   995 => x"ab4d4cc0",
   996 => x"87e8c004",
   997 => x"1ecff6c0",
   998 => x"c4029d75",
   999 => x"c24ac087",
  1000 => x"724ac187",
  1001 => x"87d6ec49",
  1002 => x"7e7086c4",
  1003 => x"056e84c1",
  1004 => x"4c7387c2",
  1005 => x"ac7385c1",
  1006 => x"87d8ff06",
  1007 => x"fe26486e",
  1008 => x"5e0e87f9",
  1009 => x"710e5c5b",
  1010 => x"0266cc4b",
  1011 => x"c04c87d8",
  1012 => x"d8028cf0",
  1013 => x"c14a7487",
  1014 => x"87d1028a",
  1015 => x"87cd028a",
  1016 => x"87c9028a",
  1017 => x"497387d9",
  1018 => x"d287c4f9",
  1019 => x"c01e7487",
  1020 => x"d4d9c149",
  1021 => x"731e7487",
  1022 => x"ccd9c149",
  1023 => x"fd86c887",
  1024 => x"5e0e87fb",
  1025 => x"0e5d5c5b",
  1026 => x"494c711e",
  1027 => x"eac291de",
  1028 => x"85714dec",
  1029 => x"c1026d97",
  1030 => x"eac287dc",
  1031 => x"7449bfd8",
  1032 => x"defd7181",
  1033 => x"487e7087",
  1034 => x"f2c00298",
  1035 => x"e0eac287",
  1036 => x"cb4a704b",
  1037 => x"eec1ff49",
  1038 => x"cb4b7487",
  1039 => x"d4e3c193",
  1040 => x"c183c483",
  1041 => x"747bfac1",
  1042 => x"e4c0c149",
  1043 => x"c17b7587",
  1044 => x"bf97c1e3",
  1045 => x"eac21e49",
  1046 => x"e5fd49e0",
  1047 => x"7486c487",
  1048 => x"ccc0c149",
  1049 => x"c149c087",
  1050 => x"c287ebc1",
  1051 => x"c048c0ea",
  1052 => x"de49c178",
  1053 => x"fc2687ca",
  1054 => x"6f4c87c1",
  1055 => x"6e696461",
  1056 => x"2e2e2e67",
  1057 => x"1e731e00",
  1058 => x"c2494a71",
  1059 => x"81bfd8ea",
  1060 => x"87effb71",
  1061 => x"029b4b70",
  1062 => x"e74987c4",
  1063 => x"eac287e9",
  1064 => x"78c048d8",
  1065 => x"d7dd49c1",
  1066 => x"87d3fb87",
  1067 => x"c149c01e",
  1068 => x"2687e3c0",
  1069 => x"4a711e4f",
  1070 => x"c191cb49",
  1071 => x"c881d4e3",
  1072 => x"c2481181",
  1073 => x"c258c4ea",
  1074 => x"c048d8ea",
  1075 => x"dc49c178",
  1076 => x"4f2687ee",
  1077 => x"0299711e",
  1078 => x"e4c187d2",
  1079 => x"50c048e9",
  1080 => x"c2c180f7",
  1081 => x"e3c140f5",
  1082 => x"87ce78cd",
  1083 => x"48e5e4c1",
  1084 => x"78c6e3c1",
  1085 => x"c2c180fc",
  1086 => x"4f2678ec",
  1087 => x"5c5b5e0e",
  1088 => x"86f40e5d",
  1089 => x"4dceddc2",
  1090 => x"a6c44cc0",
  1091 => x"c278c048",
  1092 => x"48bfd8ea",
  1093 => x"c106a8c0",
  1094 => x"ddc287c0",
  1095 => x"029848ce",
  1096 => x"c087f7c0",
  1097 => x"c81ecff6",
  1098 => x"87c70266",
  1099 => x"c048a6c4",
  1100 => x"c487c578",
  1101 => x"78c148a6",
  1102 => x"e64966c4",
  1103 => x"86c487c0",
  1104 => x"84c14d70",
  1105 => x"c14866c4",
  1106 => x"58a6c880",
  1107 => x"bfd8eac2",
  1108 => x"87c603ac",
  1109 => x"ff059d75",
  1110 => x"4cc087c9",
  1111 => x"c3029d75",
  1112 => x"f6c087dc",
  1113 => x"66c81ecf",
  1114 => x"cc87c702",
  1115 => x"78c048a6",
  1116 => x"a6cc87c5",
  1117 => x"cc78c148",
  1118 => x"c1e54966",
  1119 => x"7086c487",
  1120 => x"0298487e",
  1121 => x"4987e4c2",
  1122 => x"699781cb",
  1123 => x"0299d049",
  1124 => x"7487d4c1",
  1125 => x"c191cb49",
  1126 => x"c181d4e3",
  1127 => x"c879c5c2",
  1128 => x"51ffc381",
  1129 => x"91de4974",
  1130 => x"4deceac2",
  1131 => x"c1c28571",
  1132 => x"a5c17d97",
  1133 => x"51e0c049",
  1134 => x"97dee5c2",
  1135 => x"87d202bf",
  1136 => x"a5c284c1",
  1137 => x"dee5c24b",
  1138 => x"fe49db4a",
  1139 => x"c187d8fb",
  1140 => x"a5cd87d9",
  1141 => x"c151c049",
  1142 => x"4ba5c284",
  1143 => x"49cb4a6e",
  1144 => x"87c3fbfe",
  1145 => x"7487c4c1",
  1146 => x"c191cb49",
  1147 => x"c181d4e3",
  1148 => x"c279c2c0",
  1149 => x"bf97dee5",
  1150 => x"7487d802",
  1151 => x"c191de49",
  1152 => x"eceac284",
  1153 => x"c283714b",
  1154 => x"dd4adee5",
  1155 => x"d6fafe49",
  1156 => x"7487d887",
  1157 => x"c293de4b",
  1158 => x"cb83ecea",
  1159 => x"51c049a3",
  1160 => x"6e7384c1",
  1161 => x"fe49cb4a",
  1162 => x"c487fcf9",
  1163 => x"80c14866",
  1164 => x"c758a6c8",
  1165 => x"c5c003ac",
  1166 => x"fc056e87",
  1167 => x"487487e4",
  1168 => x"f6f48ef4",
  1169 => x"1e731e87",
  1170 => x"cb494b71",
  1171 => x"d4e3c191",
  1172 => x"4aa1c881",
  1173 => x"48c0e3c1",
  1174 => x"a1c95012",
  1175 => x"eef8c04a",
  1176 => x"ca501248",
  1177 => x"c1e3c181",
  1178 => x"c1501148",
  1179 => x"bf97c1e3",
  1180 => x"49c01e49",
  1181 => x"c287cbf5",
  1182 => x"de48c0ea",
  1183 => x"d549c178",
  1184 => x"f32687fe",
  1185 => x"5e0e87f9",
  1186 => x"0e5d5c5b",
  1187 => x"4d7186f4",
  1188 => x"c191cb49",
  1189 => x"c881d4e3",
  1190 => x"a1ca4aa1",
  1191 => x"48a6c47e",
  1192 => x"bfc8eec2",
  1193 => x"bf976e78",
  1194 => x"4c66c44b",
  1195 => x"48122c73",
  1196 => x"7058a6cc",
  1197 => x"c984c19c",
  1198 => x"49699781",
  1199 => x"c204acb7",
  1200 => x"6e4cc087",
  1201 => x"c84abf97",
  1202 => x"31724966",
  1203 => x"66c4b9ff",
  1204 => x"72487499",
  1205 => x"484a7030",
  1206 => x"eec2b071",
  1207 => x"e4c058cc",
  1208 => x"49c087cf",
  1209 => x"7587d9d4",
  1210 => x"c4f6c049",
  1211 => x"f28ef487",
  1212 => x"731e87c9",
  1213 => x"494b711e",
  1214 => x"7387cbfe",
  1215 => x"87c6fe49",
  1216 => x"1e87fcf1",
  1217 => x"4b711e73",
  1218 => x"024aa3c6",
  1219 => x"c187e3c0",
  1220 => x"87d6028a",
  1221 => x"e8c1028a",
  1222 => x"c1028a87",
  1223 => x"028a87ca",
  1224 => x"8a87efc0",
  1225 => x"c187d902",
  1226 => x"49c787e9",
  1227 => x"c187c6f6",
  1228 => x"eac287ec",
  1229 => x"78df48c0",
  1230 => x"c3d349c1",
  1231 => x"87dec187",
  1232 => x"bfd8eac2",
  1233 => x"87cbc102",
  1234 => x"c288c148",
  1235 => x"c158dcea",
  1236 => x"eac287c1",
  1237 => x"c002bfdc",
  1238 => x"eac287f9",
  1239 => x"c148bfd8",
  1240 => x"dceac280",
  1241 => x"87ebc058",
  1242 => x"bfd8eac2",
  1243 => x"c289c649",
  1244 => x"c059dcea",
  1245 => x"da03a9b7",
  1246 => x"d8eac287",
  1247 => x"d278c048",
  1248 => x"dceac287",
  1249 => x"87cb02bf",
  1250 => x"bfd8eac2",
  1251 => x"c280c648",
  1252 => x"c058dcea",
  1253 => x"87e8d149",
  1254 => x"f3c04973",
  1255 => x"deef87d3",
  1256 => x"5b5e0e87",
  1257 => x"ff0e5d5c",
  1258 => x"a6dc86d4",
  1259 => x"48a6c859",
  1260 => x"80c478c0",
  1261 => x"7866c0c1",
  1262 => x"78c180c4",
  1263 => x"78c180c4",
  1264 => x"48dceac2",
  1265 => x"eac278c1",
  1266 => x"de48bfc0",
  1267 => x"87c905a8",
  1268 => x"cc87e9f4",
  1269 => x"e6cf58a6",
  1270 => x"87e2e387",
  1271 => x"e387c4e4",
  1272 => x"4c7087d1",
  1273 => x"02acfbc0",
  1274 => x"d887fbc1",
  1275 => x"edc10566",
  1276 => x"66fcc087",
  1277 => x"6a82c44a",
  1278 => x"c11e727e",
  1279 => x"c448f4df",
  1280 => x"a1c84966",
  1281 => x"7141204a",
  1282 => x"87f905aa",
  1283 => x"4a265110",
  1284 => x"4866fcc0",
  1285 => x"78c5c9c1",
  1286 => x"81c7496a",
  1287 => x"fcc05174",
  1288 => x"81c84966",
  1289 => x"fcc051c1",
  1290 => x"81c94966",
  1291 => x"fcc051c0",
  1292 => x"81ca4966",
  1293 => x"1ec151c0",
  1294 => x"496a1ed8",
  1295 => x"f6e281c8",
  1296 => x"c186c887",
  1297 => x"c04866c0",
  1298 => x"87c701a8",
  1299 => x"c148a6c8",
  1300 => x"c187ce78",
  1301 => x"c14866c0",
  1302 => x"58a6d088",
  1303 => x"c2e287c3",
  1304 => x"48a6d087",
  1305 => x"9c7478c2",
  1306 => x"87cfcd02",
  1307 => x"c14866c8",
  1308 => x"03a866c4",
  1309 => x"dc87c4cd",
  1310 => x"78c048a6",
  1311 => x"78c080e8",
  1312 => x"7087f0e0",
  1313 => x"acd0c14c",
  1314 => x"87d7c205",
  1315 => x"e37e66c4",
  1316 => x"a6c887d4",
  1317 => x"87dbe058",
  1318 => x"ecc04c70",
  1319 => x"edc105ac",
  1320 => x"4966c887",
  1321 => x"fcc091cb",
  1322 => x"a1c48166",
  1323 => x"c84d6a4a",
  1324 => x"66c44aa1",
  1325 => x"f5c2c152",
  1326 => x"f6dfff79",
  1327 => x"9c4c7087",
  1328 => x"c087d902",
  1329 => x"d302acfb",
  1330 => x"ff557487",
  1331 => x"7087e4df",
  1332 => x"c7029c4c",
  1333 => x"acfbc087",
  1334 => x"87edff05",
  1335 => x"c255e0c0",
  1336 => x"97c055c1",
  1337 => x"4866d87d",
  1338 => x"db05a86e",
  1339 => x"4866c887",
  1340 => x"04a866cc",
  1341 => x"66c887ca",
  1342 => x"cc80c148",
  1343 => x"87c858a6",
  1344 => x"c14866cc",
  1345 => x"58a6d088",
  1346 => x"87e7deff",
  1347 => x"d0c14c70",
  1348 => x"87c805ac",
  1349 => x"c14866d4",
  1350 => x"58a6d880",
  1351 => x"02acd0c1",
  1352 => x"c487e9fd",
  1353 => x"66d84866",
  1354 => x"e0c905a8",
  1355 => x"a6e0c087",
  1356 => x"7478c048",
  1357 => x"88fbc048",
  1358 => x"98487e70",
  1359 => x"87e2c902",
  1360 => x"7088cb48",
  1361 => x"0298487e",
  1362 => x"4887cdc1",
  1363 => x"7e7088c9",
  1364 => x"c3029848",
  1365 => x"c44887fe",
  1366 => x"487e7088",
  1367 => x"87ce0298",
  1368 => x"7088c148",
  1369 => x"0298487e",
  1370 => x"c887e9c3",
  1371 => x"a6dc87d6",
  1372 => x"78f0c048",
  1373 => x"87fbdcff",
  1374 => x"ecc04c70",
  1375 => x"c4c002ac",
  1376 => x"a6e0c087",
  1377 => x"acecc05c",
  1378 => x"ff87cd02",
  1379 => x"7087e4dc",
  1380 => x"acecc04c",
  1381 => x"87f3ff05",
  1382 => x"02acecc0",
  1383 => x"ff87c4c0",
  1384 => x"c087d0dc",
  1385 => x"d01eca1e",
  1386 => x"91cb4966",
  1387 => x"4866c4c1",
  1388 => x"a6cc8071",
  1389 => x"4866c858",
  1390 => x"a6d080c4",
  1391 => x"bf66cc58",
  1392 => x"f2dcff49",
  1393 => x"de1ec187",
  1394 => x"bf66d41e",
  1395 => x"e6dcff49",
  1396 => x"7086d087",
  1397 => x"08c04849",
  1398 => x"a6e8c088",
  1399 => x"06a8c058",
  1400 => x"c087eec0",
  1401 => x"dd4866e4",
  1402 => x"e4c003a8",
  1403 => x"bf66c487",
  1404 => x"66e4c049",
  1405 => x"51e0c081",
  1406 => x"4966e4c0",
  1407 => x"66c481c1",
  1408 => x"c1c281bf",
  1409 => x"66e4c051",
  1410 => x"c481c249",
  1411 => x"c081bf66",
  1412 => x"c1486e51",
  1413 => x"6e78c5c9",
  1414 => x"d081c849",
  1415 => x"496e5166",
  1416 => x"66d481c9",
  1417 => x"ca496e51",
  1418 => x"5166dc81",
  1419 => x"c14866d0",
  1420 => x"58a6d480",
  1421 => x"cc4866c8",
  1422 => x"c004a866",
  1423 => x"66c887cb",
  1424 => x"cc80c148",
  1425 => x"d9c558a6",
  1426 => x"4866cc87",
  1427 => x"a6d088c1",
  1428 => x"87cec558",
  1429 => x"87cedcff",
  1430 => x"58a6e8c0",
  1431 => x"87c6dcff",
  1432 => x"58a6e0c0",
  1433 => x"05a8ecc0",
  1434 => x"dc87cac0",
  1435 => x"e4c048a6",
  1436 => x"c4c07866",
  1437 => x"fad8ff87",
  1438 => x"4966c887",
  1439 => x"fcc091cb",
  1440 => x"80714866",
  1441 => x"c84a7e70",
  1442 => x"ca496e82",
  1443 => x"66e4c081",
  1444 => x"4966dc51",
  1445 => x"e4c081c1",
  1446 => x"48c18966",
  1447 => x"49703071",
  1448 => x"977189c1",
  1449 => x"c8eec27a",
  1450 => x"e4c049bf",
  1451 => x"6a972966",
  1452 => x"9871484a",
  1453 => x"58a6ecc0",
  1454 => x"81c4496e",
  1455 => x"66d84d69",
  1456 => x"a866c448",
  1457 => x"87c8c002",
  1458 => x"c048a6c4",
  1459 => x"87c5c078",
  1460 => x"c148a6c4",
  1461 => x"1e66c478",
  1462 => x"751ee0c0",
  1463 => x"d6d8ff49",
  1464 => x"7086c887",
  1465 => x"acb7c04c",
  1466 => x"87d4c106",
  1467 => x"e0c08574",
  1468 => x"75897449",
  1469 => x"fddfc14b",
  1470 => x"e6fe714a",
  1471 => x"85c287e9",
  1472 => x"4866e0c0",
  1473 => x"e4c080c1",
  1474 => x"e8c058a6",
  1475 => x"81c14966",
  1476 => x"c002a970",
  1477 => x"a6c487c8",
  1478 => x"c078c048",
  1479 => x"a6c487c5",
  1480 => x"c478c148",
  1481 => x"a4c21e66",
  1482 => x"48e0c049",
  1483 => x"49708871",
  1484 => x"ff49751e",
  1485 => x"c887c0d7",
  1486 => x"a8b7c086",
  1487 => x"87c0ff01",
  1488 => x"0266e0c0",
  1489 => x"6e87d1c0",
  1490 => x"c081c949",
  1491 => x"6e5166e0",
  1492 => x"c6cac148",
  1493 => x"87ccc078",
  1494 => x"81c9496e",
  1495 => x"486e51c2",
  1496 => x"78f2cbc1",
  1497 => x"cc4866c8",
  1498 => x"c004a866",
  1499 => x"66c887cb",
  1500 => x"cc80c148",
  1501 => x"e9c058a6",
  1502 => x"4866cc87",
  1503 => x"a6d088c1",
  1504 => x"87dec058",
  1505 => x"87dbd5ff",
  1506 => x"d5c04c70",
  1507 => x"acc6c187",
  1508 => x"87c8c005",
  1509 => x"c14866d0",
  1510 => x"58a6d480",
  1511 => x"87c3d5ff",
  1512 => x"66d44c70",
  1513 => x"d880c148",
  1514 => x"9c7458a6",
  1515 => x"87cbc002",
  1516 => x"c14866c8",
  1517 => x"04a866c4",
  1518 => x"ff87fcf2",
  1519 => x"c887dbd4",
  1520 => x"a8c74866",
  1521 => x"87e5c003",
  1522 => x"48dceac2",
  1523 => x"66c878c0",
  1524 => x"c091cb49",
  1525 => x"c48166fc",
  1526 => x"4a6a4aa1",
  1527 => x"c87952c0",
  1528 => x"80c14866",
  1529 => x"c758a6cc",
  1530 => x"dbff04a8",
  1531 => x"8ed4ff87",
  1532 => x"87c7deff",
  1533 => x"64616f4c",
  1534 => x"202e2a20",
  1535 => x"00203a00",
  1536 => x"711e731e",
  1537 => x"c6029b4b",
  1538 => x"d8eac287",
  1539 => x"c778c048",
  1540 => x"d8eac21e",
  1541 => x"e3c11ebf",
  1542 => x"eac21ed4",
  1543 => x"ed49bfc0",
  1544 => x"86cc87ff",
  1545 => x"bfc0eac2",
  1546 => x"87e8e249",
  1547 => x"c8029b73",
  1548 => x"d4e3c187",
  1549 => x"cae2c049",
  1550 => x"c2ddff87",
  1551 => x"cac71e87",
  1552 => x"fe49c187",
  1553 => x"eac287fa",
  1554 => x"50c048e0",
  1555 => x"87c7eafe",
  1556 => x"cd029870",
  1557 => x"c1f3fe87",
  1558 => x"02987087",
  1559 => x"4ac187c4",
  1560 => x"4ac087c2",
  1561 => x"ce059a72",
  1562 => x"c11ec087",
  1563 => x"c049eae2",
  1564 => x"c487fbef",
  1565 => x"c287fe86",
  1566 => x"c048d8ea",
  1567 => x"c0eac278",
  1568 => x"1e78c048",
  1569 => x"49f5e2c1",
  1570 => x"87e2efc0",
  1571 => x"f8c01ec0",
  1572 => x"497087f4",
  1573 => x"87d6efc0",
  1574 => x"edc286c8",
  1575 => x"dfe2c087",
  1576 => x"d4f3c087",
  1577 => x"87f5ff87",
  1578 => x"44534f26",
  1579 => x"69616620",
  1580 => x"2e64656c",
  1581 => x"6f6f4200",
  1582 => x"676e6974",
  1583 => x"002e2e2e",
  1584 => x"00010000",
  1585 => x"20800000",
  1586 => x"74697845",
  1587 => x"42208000",
  1588 => x"006b6361",
  1589 => x"00001002",
  1590 => x"00002aac",
  1591 => x"02000000",
  1592 => x"ca000010",
  1593 => x"0000002a",
  1594 => x"10020000",
  1595 => x"2ae80000",
  1596 => x"00000000",
  1597 => x"00100200",
  1598 => x"002b0600",
  1599 => x"00000000",
  1600 => x"00001002",
  1601 => x"00002b24",
  1602 => x"02000000",
  1603 => x"42000010",
  1604 => x"0000002b",
  1605 => x"10020000",
  1606 => x"2b600000",
  1607 => x"00000000",
  1608 => x"0010b500",
  1609 => x"00000000",
  1610 => x"00000000",
  1611 => x"00001303",
  1612 => x"00000000",
  1613 => x"1e000000",
  1614 => x"c048f0fe",
  1615 => x"7909cd78",
  1616 => x"1e4f2609",
  1617 => x"48bff0fe",
  1618 => x"fe1e4f26",
  1619 => x"78c148f0",
  1620 => x"fe1e4f26",
  1621 => x"78c048f0",
  1622 => x"711e4f26",
  1623 => x"5152c04a",
  1624 => x"5e0e4f26",
  1625 => x"0e5d5c5b",
  1626 => x"4d7186f4",
  1627 => x"c17e6d97",
  1628 => x"6c974ca5",
  1629 => x"58a6c848",
  1630 => x"66c4486e",
  1631 => x"87c505a8",
  1632 => x"e6c048ff",
  1633 => x"87caff87",
  1634 => x"9749a5c2",
  1635 => x"a3714b6c",
  1636 => x"4b6b974b",
  1637 => x"6e7e6c97",
  1638 => x"c880c148",
  1639 => x"98c758a6",
  1640 => x"7058a6cc",
  1641 => x"e1fe7c97",
  1642 => x"f4487387",
  1643 => x"264d268e",
  1644 => x"264b264c",
  1645 => x"5b5e0e4f",
  1646 => x"86f40e5c",
  1647 => x"66d84c71",
  1648 => x"9affc34a",
  1649 => x"974ba4c2",
  1650 => x"a173496c",
  1651 => x"97517249",
  1652 => x"486e7e6c",
  1653 => x"a6c880c1",
  1654 => x"cc98c758",
  1655 => x"547058a6",
  1656 => x"caff8ef4",
  1657 => x"fd1e1e87",
  1658 => x"bfe087e8",
  1659 => x"e0c0494a",
  1660 => x"cb0299c0",
  1661 => x"c21e7287",
  1662 => x"fe49feed",
  1663 => x"86c487f7",
  1664 => x"7087c0fd",
  1665 => x"87c2fd7e",
  1666 => x"1e4f2626",
  1667 => x"49feedc2",
  1668 => x"c187c7fd",
  1669 => x"fc49e5e7",
  1670 => x"eec387dd",
  1671 => x"0e4f2687",
  1672 => x"5d5c5b5e",
  1673 => x"c24d710e",
  1674 => x"fc49feed",
  1675 => x"4b7087f4",
  1676 => x"04abb7c0",
  1677 => x"c387c2c3",
  1678 => x"c905abf0",
  1679 => x"c3ecc187",
  1680 => x"c278c148",
  1681 => x"e0c387e3",
  1682 => x"87c905ab",
  1683 => x"48c7ecc1",
  1684 => x"d4c278c1",
  1685 => x"c7ecc187",
  1686 => x"87c602bf",
  1687 => x"4ca3c0c2",
  1688 => x"4c7387c2",
  1689 => x"bfc3ecc1",
  1690 => x"87e0c002",
  1691 => x"b7c44974",
  1692 => x"edc19129",
  1693 => x"4a7481da",
  1694 => x"92c29acf",
  1695 => x"307248c1",
  1696 => x"baff4a70",
  1697 => x"98694872",
  1698 => x"87db7970",
  1699 => x"b7c44974",
  1700 => x"edc19129",
  1701 => x"4a7481da",
  1702 => x"92c29acf",
  1703 => x"307248c3",
  1704 => x"69484a70",
  1705 => x"757970b0",
  1706 => x"f0c0059d",
  1707 => x"48d0ff87",
  1708 => x"ff78e1c8",
  1709 => x"78c548d4",
  1710 => x"bfc7ecc1",
  1711 => x"c387c302",
  1712 => x"ecc178e0",
  1713 => x"c602bfc3",
  1714 => x"48d4ff87",
  1715 => x"ff78f0c3",
  1716 => x"0b7b0bd4",
  1717 => x"c848d0ff",
  1718 => x"e0c078e1",
  1719 => x"c7ecc178",
  1720 => x"c178c048",
  1721 => x"c048c3ec",
  1722 => x"feedc278",
  1723 => x"87f2f949",
  1724 => x"b7c04b70",
  1725 => x"fefc03ab",
  1726 => x"2648c087",
  1727 => x"264c264d",
  1728 => x"004f264b",
  1729 => x"00000000",
  1730 => x"1e000000",
  1731 => x"49724ac0",
  1732 => x"edc191c4",
  1733 => x"79c081da",
  1734 => x"b7d082c1",
  1735 => x"87ee04aa",
  1736 => x"5e0e4f26",
  1737 => x"0e5d5c5b",
  1738 => x"e5f84d71",
  1739 => x"c44a7587",
  1740 => x"c1922ab7",
  1741 => x"7582daed",
  1742 => x"c29ccf4c",
  1743 => x"4b496a94",
  1744 => x"9bc32b74",
  1745 => x"307448c2",
  1746 => x"bcff4c70",
  1747 => x"98714874",
  1748 => x"f5f77a70",
  1749 => x"fe487387",
  1750 => x"000087e1",
  1751 => x"00000000",
  1752 => x"00000000",
  1753 => x"00000000",
  1754 => x"00000000",
  1755 => x"00000000",
  1756 => x"00000000",
  1757 => x"00000000",
  1758 => x"00000000",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"ff1e0000",
  1767 => x"e1c848d0",
  1768 => x"ff487178",
  1769 => x"267808d4",
  1770 => x"d0ff1e4f",
  1771 => x"78e1c848",
  1772 => x"d4ff4871",
  1773 => x"66c47808",
  1774 => x"08d4ff48",
  1775 => x"1e4f2678",
  1776 => x"66c44a71",
  1777 => x"49721e49",
  1778 => x"ff87deff",
  1779 => x"e0c048d0",
  1780 => x"4f262678",
  1781 => x"711e731e",
  1782 => x"4966c84b",
  1783 => x"c14a731e",
  1784 => x"ff49a2e0",
  1785 => x"c42687d9",
  1786 => x"264d2687",
  1787 => x"264b264c",
  1788 => x"d4ff1e4f",
  1789 => x"7affc34a",
  1790 => x"c048d0ff",
  1791 => x"7ade78e1",
  1792 => x"bfc8eec2",
  1793 => x"c848497a",
  1794 => x"717a7028",
  1795 => x"7028d048",
  1796 => x"d848717a",
  1797 => x"ff7a7028",
  1798 => x"e0c048d0",
  1799 => x"1e4f2678",
  1800 => x"c848d0ff",
  1801 => x"487178c9",
  1802 => x"7808d4ff",
  1803 => x"711e4f26",
  1804 => x"87eb494a",
  1805 => x"c848d0ff",
  1806 => x"1e4f2678",
  1807 => x"4b711e73",
  1808 => x"bfd8eec2",
  1809 => x"c287c302",
  1810 => x"d0ff87eb",
  1811 => x"78c9c848",
  1812 => x"e0c04873",
  1813 => x"08d4ffb0",
  1814 => x"cceec278",
  1815 => x"c878c048",
  1816 => x"87c50266",
  1817 => x"c249ffc3",
  1818 => x"c249c087",
  1819 => x"cc59d4ee",
  1820 => x"87c60266",
  1821 => x"4ad5d5c5",
  1822 => x"ffcf87c4",
  1823 => x"eec24aff",
  1824 => x"eec25ad8",
  1825 => x"78c148d8",
  1826 => x"4d2687c4",
  1827 => x"4b264c26",
  1828 => x"5e0e4f26",
  1829 => x"0e5d5c5b",
  1830 => x"eec24a71",
  1831 => x"724cbfd4",
  1832 => x"87cb029a",
  1833 => x"c191c849",
  1834 => x"714bf1f0",
  1835 => x"c187c483",
  1836 => x"c04bf1f4",
  1837 => x"7449134d",
  1838 => x"d0eec299",
  1839 => x"b87148bf",
  1840 => x"7808d4ff",
  1841 => x"852cb7c1",
  1842 => x"04adb7c8",
  1843 => x"eec287e7",
  1844 => x"c848bfcc",
  1845 => x"d0eec280",
  1846 => x"87eefe58",
  1847 => x"711e731e",
  1848 => x"9a4a134b",
  1849 => x"7287cb02",
  1850 => x"87e6fe49",
  1851 => x"059a4a13",
  1852 => x"d9fe87f5",
  1853 => x"eec21e87",
  1854 => x"c249bfcc",
  1855 => x"c148ccee",
  1856 => x"c0c478a1",
  1857 => x"db03a9b7",
  1858 => x"48d4ff87",
  1859 => x"bfd0eec2",
  1860 => x"cceec278",
  1861 => x"eec249bf",
  1862 => x"a1c148cc",
  1863 => x"b7c0c478",
  1864 => x"87e504a9",
  1865 => x"c848d0ff",
  1866 => x"d8eec278",
  1867 => x"2678c048",
  1868 => x"0000004f",
  1869 => x"00000000",
  1870 => x"00000000",
  1871 => x"00005f5f",
  1872 => x"03030000",
  1873 => x"00030300",
  1874 => x"7f7f1400",
  1875 => x"147f7f14",
  1876 => x"2e240000",
  1877 => x"123a6b6b",
  1878 => x"366a4c00",
  1879 => x"32566c18",
  1880 => x"4f7e3000",
  1881 => x"683a7759",
  1882 => x"04000040",
  1883 => x"00000307",
  1884 => x"1c000000",
  1885 => x"0041633e",
  1886 => x"41000000",
  1887 => x"001c3e63",
  1888 => x"3e2a0800",
  1889 => x"2a3e1c1c",
  1890 => x"08080008",
  1891 => x"08083e3e",
  1892 => x"80000000",
  1893 => x"000060e0",
  1894 => x"08080000",
  1895 => x"08080808",
  1896 => x"00000000",
  1897 => x"00006060",
  1898 => x"30604000",
  1899 => x"03060c18",
  1900 => x"7f3e0001",
  1901 => x"3e7f4d59",
  1902 => x"06040000",
  1903 => x"00007f7f",
  1904 => x"63420000",
  1905 => x"464f5971",
  1906 => x"63220000",
  1907 => x"367f4949",
  1908 => x"161c1800",
  1909 => x"107f7f13",
  1910 => x"67270000",
  1911 => x"397d4545",
  1912 => x"7e3c0000",
  1913 => x"3079494b",
  1914 => x"01010000",
  1915 => x"070f7971",
  1916 => x"7f360000",
  1917 => x"367f4949",
  1918 => x"4f060000",
  1919 => x"1e3f6949",
  1920 => x"00000000",
  1921 => x"00006666",
  1922 => x"80000000",
  1923 => x"000066e6",
  1924 => x"08080000",
  1925 => x"22221414",
  1926 => x"14140000",
  1927 => x"14141414",
  1928 => x"22220000",
  1929 => x"08081414",
  1930 => x"03020000",
  1931 => x"060f5951",
  1932 => x"417f3e00",
  1933 => x"1e1f555d",
  1934 => x"7f7e0000",
  1935 => x"7e7f0909",
  1936 => x"7f7f0000",
  1937 => x"367f4949",
  1938 => x"3e1c0000",
  1939 => x"41414163",
  1940 => x"7f7f0000",
  1941 => x"1c3e6341",
  1942 => x"7f7f0000",
  1943 => x"41414949",
  1944 => x"7f7f0000",
  1945 => x"01010909",
  1946 => x"7f3e0000",
  1947 => x"7a7b4941",
  1948 => x"7f7f0000",
  1949 => x"7f7f0808",
  1950 => x"41000000",
  1951 => x"00417f7f",
  1952 => x"60200000",
  1953 => x"3f7f4040",
  1954 => x"087f7f00",
  1955 => x"4163361c",
  1956 => x"7f7f0000",
  1957 => x"40404040",
  1958 => x"067f7f00",
  1959 => x"7f7f060c",
  1960 => x"067f7f00",
  1961 => x"7f7f180c",
  1962 => x"7f3e0000",
  1963 => x"3e7f4141",
  1964 => x"7f7f0000",
  1965 => x"060f0909",
  1966 => x"417f3e00",
  1967 => x"407e7f61",
  1968 => x"7f7f0000",
  1969 => x"667f1909",
  1970 => x"6f260000",
  1971 => x"327b594d",
  1972 => x"01010000",
  1973 => x"01017f7f",
  1974 => x"7f3f0000",
  1975 => x"3f7f4040",
  1976 => x"3f0f0000",
  1977 => x"0f3f7070",
  1978 => x"307f7f00",
  1979 => x"7f7f3018",
  1980 => x"36634100",
  1981 => x"63361c1c",
  1982 => x"06030141",
  1983 => x"03067c7c",
  1984 => x"59716101",
  1985 => x"4143474d",
  1986 => x"7f000000",
  1987 => x"0041417f",
  1988 => x"06030100",
  1989 => x"6030180c",
  1990 => x"41000040",
  1991 => x"007f7f41",
  1992 => x"060c0800",
  1993 => x"080c0603",
  1994 => x"80808000",
  1995 => x"80808080",
  1996 => x"00000000",
  1997 => x"00040703",
  1998 => x"74200000",
  1999 => x"787c5454",
  2000 => x"7f7f0000",
  2001 => x"387c4444",
  2002 => x"7c380000",
  2003 => x"00444444",
  2004 => x"7c380000",
  2005 => x"7f7f4444",
  2006 => x"7c380000",
  2007 => x"185c5454",
  2008 => x"7e040000",
  2009 => x"0005057f",
  2010 => x"bc180000",
  2011 => x"7cfca4a4",
  2012 => x"7f7f0000",
  2013 => x"787c0404",
  2014 => x"00000000",
  2015 => x"00407d3d",
  2016 => x"80800000",
  2017 => x"007dfd80",
  2018 => x"7f7f0000",
  2019 => x"446c3810",
  2020 => x"00000000",
  2021 => x"00407f3f",
  2022 => x"0c7c7c00",
  2023 => x"787c0c18",
  2024 => x"7c7c0000",
  2025 => x"787c0404",
  2026 => x"7c380000",
  2027 => x"387c4444",
  2028 => x"fcfc0000",
  2029 => x"183c2424",
  2030 => x"3c180000",
  2031 => x"fcfc2424",
  2032 => x"7c7c0000",
  2033 => x"080c0404",
  2034 => x"5c480000",
  2035 => x"20745454",
  2036 => x"3f040000",
  2037 => x"0044447f",
  2038 => x"7c3c0000",
  2039 => x"7c7c4040",
  2040 => x"3c1c0000",
  2041 => x"1c3c6060",
  2042 => x"607c3c00",
  2043 => x"3c7c6030",
  2044 => x"386c4400",
  2045 => x"446c3810",
  2046 => x"bc1c0000",
  2047 => x"1c3c60e0",
  2048 => x"64440000",
  2049 => x"444c5c74",
  2050 => x"08080000",
  2051 => x"4141773e",
  2052 => x"00000000",
  2053 => x"00007f7f",
  2054 => x"41410000",
  2055 => x"08083e77",
  2056 => x"01010200",
  2057 => x"01020203",
  2058 => x"7f7f7f00",
  2059 => x"7f7f7f7f",
  2060 => x"1c080800",
  2061 => x"7f3e3e1c",
  2062 => x"3e7f7f7f",
  2063 => x"081c1c3e",
  2064 => x"18100008",
  2065 => x"10187c7c",
  2066 => x"30100000",
  2067 => x"10307c7c",
  2068 => x"60301000",
  2069 => x"061e7860",
  2070 => x"3c664200",
  2071 => x"42663c18",
  2072 => x"6a387800",
  2073 => x"386cc6c2",
  2074 => x"00006000",
  2075 => x"60000060",
  2076 => x"5b5e0e00",
  2077 => x"1e0e5d5c",
  2078 => x"eec24c71",
  2079 => x"c04dbfdd",
  2080 => x"741ec04b",
  2081 => x"87c702ab",
  2082 => x"c048a6c4",
  2083 => x"c487c578",
  2084 => x"78c148a6",
  2085 => x"731e66c4",
  2086 => x"87dfee49",
  2087 => x"e0c086c8",
  2088 => x"87eeef49",
  2089 => x"6a4aa5c4",
  2090 => x"87f0f049",
  2091 => x"cb87c6f1",
  2092 => x"c883c185",
  2093 => x"ff04abb7",
  2094 => x"262687c7",
  2095 => x"264c264d",
  2096 => x"1e4f264b",
  2097 => x"eec24a71",
  2098 => x"eec25ae1",
  2099 => x"78c748e1",
  2100 => x"87ddfe49",
  2101 => x"731e4f26",
  2102 => x"c04a711e",
  2103 => x"d303aab7",
  2104 => x"d8d3c287",
  2105 => x"87c405bf",
  2106 => x"87c24bc1",
  2107 => x"d3c24bc0",
  2108 => x"87c45bdc",
  2109 => x"5adcd3c2",
  2110 => x"bfd8d3c2",
  2111 => x"c19ac14a",
  2112 => x"ec49a2c0",
  2113 => x"48fc87e8",
  2114 => x"bfd8d3c2",
  2115 => x"87effe78",
  2116 => x"c44a711e",
  2117 => x"49721e66",
  2118 => x"2687f9ea",
  2119 => x"ff1e4f26",
  2120 => x"ffc348d4",
  2121 => x"48d0ff78",
  2122 => x"ff78e1c0",
  2123 => x"78c148d4",
  2124 => x"30c44871",
  2125 => x"7808d4ff",
  2126 => x"c048d0ff",
  2127 => x"4f2678e0",
  2128 => x"5c5b5e0e",
  2129 => x"86f40e5d",
  2130 => x"c048a6c4",
  2131 => x"bfec4b78",
  2132 => x"ddeec27e",
  2133 => x"bfe84dbf",
  2134 => x"d8d3c24c",
  2135 => x"fee249bf",
  2136 => x"49eecb87",
  2137 => x"cc87f9cd",
  2138 => x"49c758a6",
  2139 => x"7087f3e6",
  2140 => x"87c80598",
  2141 => x"99c1496e",
  2142 => x"87c3c102",
  2143 => x"bfec4bc1",
  2144 => x"d8d3c27e",
  2145 => x"d6e249bf",
  2146 => x"4966c887",
  2147 => x"7087ddcd",
  2148 => x"87d80298",
  2149 => x"bfc0d3c2",
  2150 => x"c2b9c149",
  2151 => x"7159c4d3",
  2152 => x"cb87fbfd",
  2153 => x"f7cc49ee",
  2154 => x"58a6cc87",
  2155 => x"f1e549c7",
  2156 => x"05987087",
  2157 => x"6e87c5ff",
  2158 => x"0599c149",
  2159 => x"7387fdfe",
  2160 => x"87d0029b",
  2161 => x"cdfc49ff",
  2162 => x"49dac187",
  2163 => x"c487d3e5",
  2164 => x"78c148a6",
  2165 => x"bfd8d3c2",
  2166 => x"87d9c105",
  2167 => x"c848a6c4",
  2168 => x"c278c0c0",
  2169 => x"6e7ec4d3",
  2170 => x"6e49bf97",
  2171 => x"7080c148",
  2172 => x"ede4717e",
  2173 => x"02987087",
  2174 => x"66c487c3",
  2175 => x"4866c4b4",
  2176 => x"c828b7c1",
  2177 => x"987058a6",
  2178 => x"87dbff05",
  2179 => x"e449fdc3",
  2180 => x"fac387d0",
  2181 => x"87cae449",
  2182 => x"ffc34974",
  2183 => x"c01e7199",
  2184 => x"87ecfb49",
  2185 => x"b7c84974",
  2186 => x"c11e7129",
  2187 => x"87e0fb49",
  2188 => x"f4c886c8",
  2189 => x"c3497487",
  2190 => x"b7c899ff",
  2191 => x"74b4712c",
  2192 => x"87df029c",
  2193 => x"bfd4d3c2",
  2194 => x"87e0ca49",
  2195 => x"c0059870",
  2196 => x"4cc087c4",
  2197 => x"e0c287d3",
  2198 => x"87c4ca49",
  2199 => x"58d8d3c2",
  2200 => x"c287c6c0",
  2201 => x"c048d4d3",
  2202 => x"c2497478",
  2203 => x"cec00599",
  2204 => x"49ebc387",
  2205 => x"7087ebe2",
  2206 => x"0299c249",
  2207 => x"c187cfc0",
  2208 => x"6e7ea5d8",
  2209 => x"c5c002bf",
  2210 => x"49fb4b87",
  2211 => x"49740f73",
  2212 => x"c00599c1",
  2213 => x"f4c387ce",
  2214 => x"87c6e249",
  2215 => x"99c24970",
  2216 => x"87cfc002",
  2217 => x"7ea5d8c1",
  2218 => x"c002bf6e",
  2219 => x"fa4b87c5",
  2220 => x"740f7349",
  2221 => x"0599c849",
  2222 => x"c387cec0",
  2223 => x"e1e149f5",
  2224 => x"c2497087",
  2225 => x"e5c00299",
  2226 => x"e1eec287",
  2227 => x"cac002bf",
  2228 => x"88c14887",
  2229 => x"58e5eec2",
  2230 => x"c187cec0",
  2231 => x"6a4aa5d8",
  2232 => x"87c5c002",
  2233 => x"7349ff4b",
  2234 => x"48a6c40f",
  2235 => x"497478c1",
  2236 => x"c00599c4",
  2237 => x"f2c387ce",
  2238 => x"87e6e049",
  2239 => x"99c24970",
  2240 => x"87ecc002",
  2241 => x"bfe1eec2",
  2242 => x"b7c7487e",
  2243 => x"cbc003a8",
  2244 => x"c1486e87",
  2245 => x"e5eec280",
  2246 => x"87cfc058",
  2247 => x"7ea5d8c1",
  2248 => x"c002bf6e",
  2249 => x"fe4b87c5",
  2250 => x"c40f7349",
  2251 => x"78c148a6",
  2252 => x"ff49fdc3",
  2253 => x"7087ebdf",
  2254 => x"0299c249",
  2255 => x"c287e5c0",
  2256 => x"02bfe1ee",
  2257 => x"c287c9c0",
  2258 => x"c048e1ee",
  2259 => x"87cfc078",
  2260 => x"7ea5d8c1",
  2261 => x"c002bf6e",
  2262 => x"fd4b87c5",
  2263 => x"c40f7349",
  2264 => x"78c148a6",
  2265 => x"ff49fac3",
  2266 => x"7087f7de",
  2267 => x"0299c249",
  2268 => x"c287e9c0",
  2269 => x"48bfe1ee",
  2270 => x"03a8b7c7",
  2271 => x"c287c9c0",
  2272 => x"c748e1ee",
  2273 => x"87cfc078",
  2274 => x"7ea5d8c1",
  2275 => x"c002bf6e",
  2276 => x"fc4b87c5",
  2277 => x"c40f7349",
  2278 => x"78c148a6",
  2279 => x"eec24bc0",
  2280 => x"50c048dc",
  2281 => x"c449eecb",
  2282 => x"a6cc87f6",
  2283 => x"dceec258",
  2284 => x"c105bf97",
  2285 => x"497487de",
  2286 => x"0599f0c3",
  2287 => x"c187cdc0",
  2288 => x"ddff49da",
  2289 => x"987087dc",
  2290 => x"87c8c102",
  2291 => x"bfe84bc1",
  2292 => x"ffc3494c",
  2293 => x"2cb7c899",
  2294 => x"d3c2b471",
  2295 => x"ff49bfd8",
  2296 => x"c887fcd8",
  2297 => x"c3c44966",
  2298 => x"02987087",
  2299 => x"c287c6c0",
  2300 => x"c148dcee",
  2301 => x"dceec250",
  2302 => x"c005bf97",
  2303 => x"497487d6",
  2304 => x"0599f0c3",
  2305 => x"c187c5ff",
  2306 => x"dcff49da",
  2307 => x"987087d4",
  2308 => x"87f8fe05",
  2309 => x"c0029b73",
  2310 => x"a6c887dc",
  2311 => x"e1eec248",
  2312 => x"66c878bf",
  2313 => x"7591cb49",
  2314 => x"bf6e7ea1",
  2315 => x"87c6c002",
  2316 => x"4966c84b",
  2317 => x"66c40f73",
  2318 => x"87c8c002",
  2319 => x"bfe1eec2",
  2320 => x"87edf049",
  2321 => x"bfdcd3c2",
  2322 => x"87ddc002",
  2323 => x"87dcc249",
  2324 => x"c0029870",
  2325 => x"eec287d3",
  2326 => x"f049bfe1",
  2327 => x"49c087d3",
  2328 => x"c287f3f1",
  2329 => x"c048dcd3",
  2330 => x"f18ef478",
  2331 => x"5e0e87cd",
  2332 => x"0e5d5c5b",
  2333 => x"c24c711e",
  2334 => x"49bfddee",
  2335 => x"4da1cdc1",
  2336 => x"6981d1c1",
  2337 => x"029c747e",
  2338 => x"a5c487cf",
  2339 => x"c27b744b",
  2340 => x"49bfddee",
  2341 => x"6e87ecf0",
  2342 => x"059c747b",
  2343 => x"4bc087c4",
  2344 => x"4bc187c2",
  2345 => x"edf04973",
  2346 => x"0266d487",
  2347 => x"c04987c8",
  2348 => x"4a7087ee",
  2349 => x"4ac087c2",
  2350 => x"5ae0d3c2",
  2351 => x"87fbef26",
  2352 => x"00000000",
  2353 => x"14111258",
  2354 => x"231c1b1d",
  2355 => x"9491595a",
  2356 => x"f4ebf2f5",
  2357 => x"00000000",
  2358 => x"00000000",
  2359 => x"00000000",
  2360 => x"ff4a711e",
  2361 => x"7249bfc8",
  2362 => x"4f2648a1",
  2363 => x"bfc8ff1e",
  2364 => x"c0c0fe89",
  2365 => x"a9c0c0c0",
  2366 => x"c087c401",
  2367 => x"c187c24a",
  2368 => x"2648724a",
  2369 => x"5b5e0e4f",
  2370 => x"710e5d5c",
  2371 => x"4cd4ff4b",
  2372 => x"c04866d0",
  2373 => x"ff49d678",
  2374 => x"c387ffd9",
  2375 => x"496c7cff",
  2376 => x"7199ffc3",
  2377 => x"f0c3494d",
  2378 => x"a9e0c199",
  2379 => x"c387cb05",
  2380 => x"486c7cff",
  2381 => x"66d098c3",
  2382 => x"ffc37808",
  2383 => x"494a6c7c",
  2384 => x"ffc331c8",
  2385 => x"714a6c7c",
  2386 => x"c84972b2",
  2387 => x"7cffc331",
  2388 => x"b2714a6c",
  2389 => x"31c84972",
  2390 => x"6c7cffc3",
  2391 => x"ffb2714a",
  2392 => x"e0c048d0",
  2393 => x"029b7378",
  2394 => x"7b7287c2",
  2395 => x"4d264875",
  2396 => x"4b264c26",
  2397 => x"261e4f26",
  2398 => x"5b5e0e4f",
  2399 => x"86f80e5c",
  2400 => x"a6c81e76",
  2401 => x"87fdfd49",
  2402 => x"4b7086c4",
  2403 => x"a8c2486e",
  2404 => x"87f0c203",
  2405 => x"f0c34a73",
  2406 => x"aad0c19a",
  2407 => x"c187c702",
  2408 => x"c205aae0",
  2409 => x"497387de",
  2410 => x"c30299c8",
  2411 => x"87c6ff87",
  2412 => x"9cc34c73",
  2413 => x"c105acc2",
  2414 => x"66c487c2",
  2415 => x"7131c949",
  2416 => x"4a66c41e",
  2417 => x"eec292d4",
  2418 => x"817249e5",
  2419 => x"87f7cffe",
  2420 => x"d7ff49d8",
  2421 => x"c0c887c4",
  2422 => x"ceddc21e",
  2423 => x"fdebfd49",
  2424 => x"48d0ff87",
  2425 => x"c278e0c0",
  2426 => x"cc1ecedd",
  2427 => x"92d44a66",
  2428 => x"49e5eec2",
  2429 => x"cdfe8172",
  2430 => x"86cc87ff",
  2431 => x"c105acc1",
  2432 => x"66c487c2",
  2433 => x"7131c949",
  2434 => x"4a66c41e",
  2435 => x"eec292d4",
  2436 => x"817249e5",
  2437 => x"87efcefe",
  2438 => x"1eceddc2",
  2439 => x"d44a66c8",
  2440 => x"e5eec292",
  2441 => x"fe817249",
  2442 => x"d787c0cc",
  2443 => x"e9d5ff49",
  2444 => x"1ec0c887",
  2445 => x"49ceddc2",
  2446 => x"87fbe9fd",
  2447 => x"d0ff86cc",
  2448 => x"78e0c048",
  2449 => x"e7fc8ef8",
  2450 => x"5b5e0e87",
  2451 => x"710e5d5c",
  2452 => x"4cd4ff4a",
  2453 => x"c34d66d0",
  2454 => x"c506adb7",
  2455 => x"c148c087",
  2456 => x"1e7287e1",
  2457 => x"93d44b75",
  2458 => x"83e5eec2",
  2459 => x"c6fe4973",
  2460 => x"83c887c7",
  2461 => x"d0ff4b6b",
  2462 => x"78e1c848",
  2463 => x"48737cdd",
  2464 => x"7098ffc3",
  2465 => x"c849737c",
  2466 => x"487129b7",
  2467 => x"7098ffc3",
  2468 => x"d049737c",
  2469 => x"487129b7",
  2470 => x"7098ffc3",
  2471 => x"d848737c",
  2472 => x"7c7028b7",
  2473 => x"7c7c7cc0",
  2474 => x"7c7c7c7c",
  2475 => x"7c7c7c7c",
  2476 => x"48d0ff7c",
  2477 => x"7578e0c0",
  2478 => x"ff49dc1e",
  2479 => x"c887c0d4",
  2480 => x"fa487386",
  2481 => x"731e87e8",
  2482 => x"1e4bc01e",
  2483 => x"bfc7dcc2",
  2484 => x"87f5fd49",
  2485 => x"dcc286c4",
  2486 => x"fe49bfcb",
  2487 => x"7087d0dd",
  2488 => x"87c40598",
  2489 => x"4bf4dbc2",
  2490 => x"87c44873",
  2491 => x"4c264d26",
  2492 => x"4f264b26",
  2493 => x"204d4f52",
  2494 => x"64616f6c",
  2495 => x"20676e69",
  2496 => x"6c696166",
  2497 => x"0f006465",
  2498 => x"1b000027",
  2499 => x"42000027",
  2500 => x"20204342",
  2501 => x"56202020",
  2502 => x"42004448",
  2503 => x"20204342",
  2504 => x"52202020",
  2505 => x"52004d4f",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
