
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d0",x"ef",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"d0",x"ef",x"c2"),
    14 => (x"48",x"e8",x"dc",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"f2",x"df"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"48",x"72"),
    82 => (x"c2",x"7c",x"70",x"98"),
    83 => (x"05",x"bf",x"e8",x"dc"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"71",x"29",x"d8",x"49"),
    88 => (x"98",x"ff",x"c3",x"48"),
    89 => (x"66",x"d0",x"7c",x"70"),
    90 => (x"71",x"29",x"d0",x"49"),
    91 => (x"98",x"ff",x"c3",x"48"),
    92 => (x"66",x"d0",x"7c",x"70"),
    93 => (x"71",x"29",x"c8",x"49"),
    94 => (x"98",x"ff",x"c3",x"48"),
    95 => (x"66",x"d0",x"7c",x"70"),
    96 => (x"98",x"ff",x"c3",x"48"),
    97 => (x"49",x"72",x"7c",x"70"),
    98 => (x"48",x"71",x"29",x"d0"),
    99 => (x"70",x"98",x"ff",x"c3"),
   100 => (x"c9",x"4b",x"6c",x"7c"),
   101 => (x"c3",x"4d",x"ff",x"f0"),
   102 => (x"d0",x"05",x"ab",x"ff"),
   103 => (x"7c",x"ff",x"c3",x"87"),
   104 => (x"8d",x"c1",x"4b",x"6c"),
   105 => (x"c3",x"87",x"c6",x"02"),
   106 => (x"f0",x"02",x"ab",x"ff"),
   107 => (x"fd",x"48",x"73",x"87"),
   108 => (x"c0",x"1e",x"87",x"ff"),
   109 => (x"48",x"d4",x"ff",x"49"),
   110 => (x"c1",x"78",x"ff",x"c3"),
   111 => (x"b7",x"c8",x"c3",x"81"),
   112 => (x"87",x"f1",x"04",x"a9"),
   113 => (x"73",x"1e",x"4f",x"26"),
   114 => (x"c4",x"87",x"e7",x"1e"),
   115 => (x"c0",x"4b",x"df",x"f8"),
   116 => (x"f0",x"ff",x"c0",x"1e"),
   117 => (x"fd",x"49",x"f7",x"c1"),
   118 => (x"86",x"c4",x"87",x"df"),
   119 => (x"c0",x"05",x"a8",x"c1"),
   120 => (x"d4",x"ff",x"87",x"ea"),
   121 => (x"78",x"ff",x"c3",x"48"),
   122 => (x"c0",x"c0",x"c0",x"c1"),
   123 => (x"c0",x"1e",x"c0",x"c0"),
   124 => (x"e9",x"c1",x"f0",x"e1"),
   125 => (x"87",x"c1",x"fd",x"49"),
   126 => (x"98",x"70",x"86",x"c4"),
   127 => (x"ff",x"87",x"ca",x"05"),
   128 => (x"ff",x"c3",x"48",x"d4"),
   129 => (x"cb",x"48",x"c1",x"78"),
   130 => (x"87",x"e6",x"fe",x"87"),
   131 => (x"fe",x"05",x"8b",x"c1"),
   132 => (x"48",x"c0",x"87",x"fd"),
   133 => (x"1e",x"87",x"de",x"fc"),
   134 => (x"d4",x"ff",x"1e",x"73"),
   135 => (x"78",x"ff",x"c3",x"48"),
   136 => (x"1e",x"c0",x"4b",x"d3"),
   137 => (x"c1",x"f0",x"ff",x"c0"),
   138 => (x"cc",x"fc",x"49",x"c1"),
   139 => (x"70",x"86",x"c4",x"87"),
   140 => (x"87",x"ca",x"05",x"98"),
   141 => (x"c3",x"48",x"d4",x"ff"),
   142 => (x"48",x"c1",x"78",x"ff"),
   143 => (x"f1",x"fd",x"87",x"cb"),
   144 => (x"05",x"8b",x"c1",x"87"),
   145 => (x"c0",x"87",x"db",x"ff"),
   146 => (x"87",x"e9",x"fb",x"48"),
   147 => (x"5c",x"5b",x"5e",x"0e"),
   148 => (x"4c",x"d4",x"ff",x"0e"),
   149 => (x"c6",x"87",x"db",x"fd"),
   150 => (x"e1",x"c0",x"1e",x"ea"),
   151 => (x"49",x"c8",x"c1",x"f0"),
   152 => (x"c4",x"87",x"d6",x"fb"),
   153 => (x"02",x"a8",x"c1",x"86"),
   154 => (x"ea",x"fe",x"87",x"c8"),
   155 => (x"c1",x"48",x"c0",x"87"),
   156 => (x"d2",x"fa",x"87",x"e2"),
   157 => (x"cf",x"49",x"70",x"87"),
   158 => (x"c6",x"99",x"ff",x"ff"),
   159 => (x"c8",x"02",x"a9",x"ea"),
   160 => (x"87",x"d3",x"fe",x"87"),
   161 => (x"cb",x"c1",x"48",x"c0"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"fc",x"4b",x"f1",x"c0"),
   164 => (x"98",x"70",x"87",x"f4"),
   165 => (x"87",x"eb",x"c0",x"02"),
   166 => (x"ff",x"c0",x"1e",x"c0"),
   167 => (x"49",x"fa",x"c1",x"f0"),
   168 => (x"c4",x"87",x"d6",x"fa"),
   169 => (x"05",x"98",x"70",x"86"),
   170 => (x"ff",x"c3",x"87",x"d9"),
   171 => (x"c3",x"49",x"6c",x"7c"),
   172 => (x"7c",x"7c",x"7c",x"ff"),
   173 => (x"99",x"c0",x"c1",x"7c"),
   174 => (x"c1",x"87",x"c4",x"02"),
   175 => (x"c0",x"87",x"d5",x"48"),
   176 => (x"c2",x"87",x"d1",x"48"),
   177 => (x"87",x"c4",x"05",x"ab"),
   178 => (x"87",x"c8",x"48",x"c0"),
   179 => (x"fe",x"05",x"8b",x"c1"),
   180 => (x"48",x"c0",x"87",x"fd"),
   181 => (x"1e",x"87",x"dc",x"f9"),
   182 => (x"dc",x"c2",x"1e",x"73"),
   183 => (x"78",x"c1",x"48",x"e8"),
   184 => (x"d0",x"ff",x"4b",x"c7"),
   185 => (x"fb",x"78",x"c2",x"48"),
   186 => (x"d0",x"ff",x"87",x"c8"),
   187 => (x"c0",x"78",x"c3",x"48"),
   188 => (x"d0",x"e5",x"c0",x"1e"),
   189 => (x"f8",x"49",x"c0",x"c1"),
   190 => (x"86",x"c4",x"87",x"ff"),
   191 => (x"c1",x"05",x"a8",x"c1"),
   192 => (x"ab",x"c2",x"4b",x"87"),
   193 => (x"c0",x"87",x"c5",x"05"),
   194 => (x"87",x"f9",x"c0",x"48"),
   195 => (x"ff",x"05",x"8b",x"c1"),
   196 => (x"f7",x"fc",x"87",x"d0"),
   197 => (x"ec",x"dc",x"c2",x"87"),
   198 => (x"05",x"98",x"70",x"58"),
   199 => (x"1e",x"c1",x"87",x"cd"),
   200 => (x"c1",x"f0",x"ff",x"c0"),
   201 => (x"d0",x"f8",x"49",x"d0"),
   202 => (x"ff",x"86",x"c4",x"87"),
   203 => (x"ff",x"c3",x"48",x"d4"),
   204 => (x"87",x"dd",x"c4",x"78"),
   205 => (x"58",x"f0",x"dc",x"c2"),
   206 => (x"c2",x"48",x"d0",x"ff"),
   207 => (x"48",x"d4",x"ff",x"78"),
   208 => (x"c1",x"78",x"ff",x"c3"),
   209 => (x"87",x"ed",x"f7",x"48"),
   210 => (x"5c",x"5b",x"5e",x"0e"),
   211 => (x"4a",x"71",x"0e",x"5d"),
   212 => (x"ff",x"4d",x"ff",x"c3"),
   213 => (x"7c",x"75",x"4c",x"d4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"7c",x"75",x"78",x"c3"),
   216 => (x"ff",x"c0",x"1e",x"72"),
   217 => (x"49",x"d8",x"c1",x"f0"),
   218 => (x"c4",x"87",x"ce",x"f7"),
   219 => (x"02",x"98",x"70",x"86"),
   220 => (x"48",x"c1",x"87",x"c5"),
   221 => (x"75",x"87",x"ee",x"c0"),
   222 => (x"7c",x"fe",x"c3",x"7c"),
   223 => (x"d4",x"1e",x"c0",x"c8"),
   224 => (x"f2",x"f4",x"49",x"66"),
   225 => (x"75",x"86",x"c4",x"87"),
   226 => (x"75",x"7c",x"75",x"7c"),
   227 => (x"e0",x"da",x"d8",x"7c"),
   228 => (x"6c",x"7c",x"75",x"4b"),
   229 => (x"c1",x"87",x"c5",x"05"),
   230 => (x"87",x"f5",x"05",x"8b"),
   231 => (x"d0",x"ff",x"7c",x"75"),
   232 => (x"c0",x"78",x"c2",x"48"),
   233 => (x"87",x"c9",x"f6",x"48"),
   234 => (x"5c",x"5b",x"5e",x"0e"),
   235 => (x"4b",x"71",x"0e",x"5d"),
   236 => (x"ee",x"c5",x"4c",x"c0"),
   237 => (x"ff",x"4a",x"df",x"cd"),
   238 => (x"ff",x"c3",x"48",x"d4"),
   239 => (x"c3",x"48",x"68",x"78"),
   240 => (x"c0",x"05",x"a8",x"fe"),
   241 => (x"d4",x"ff",x"87",x"fe"),
   242 => (x"02",x"9b",x"73",x"4d"),
   243 => (x"66",x"d0",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c8"),
   246 => (x"d0",x"ff",x"87",x"d6"),
   247 => (x"78",x"d1",x"c4",x"48"),
   248 => (x"d0",x"7d",x"ff",x"c3"),
   249 => (x"88",x"c1",x"48",x"66"),
   250 => (x"70",x"58",x"a6",x"d4"),
   251 => (x"87",x"f0",x"05",x"98"),
   252 => (x"c3",x"48",x"d4",x"ff"),
   253 => (x"73",x"78",x"78",x"ff"),
   254 => (x"87",x"c5",x"05",x"9b"),
   255 => (x"d0",x"48",x"d0",x"ff"),
   256 => (x"4c",x"4a",x"c1",x"78"),
   257 => (x"fe",x"05",x"8a",x"c1"),
   258 => (x"48",x"74",x"87",x"ed"),
   259 => (x"1e",x"87",x"e2",x"f4"),
   260 => (x"4a",x"71",x"1e",x"73"),
   261 => (x"d4",x"ff",x"4b",x"c0"),
   262 => (x"78",x"ff",x"c3",x"48"),
   263 => (x"c4",x"48",x"d0",x"ff"),
   264 => (x"d4",x"ff",x"78",x"c3"),
   265 => (x"78",x"ff",x"c3",x"48"),
   266 => (x"ff",x"c0",x"1e",x"72"),
   267 => (x"49",x"d1",x"c1",x"f0"),
   268 => (x"c4",x"87",x"c6",x"f4"),
   269 => (x"05",x"98",x"70",x"86"),
   270 => (x"c0",x"c8",x"87",x"d2"),
   271 => (x"49",x"66",x"cc",x"1e"),
   272 => (x"c4",x"87",x"e5",x"fd"),
   273 => (x"ff",x"4b",x"70",x"86"),
   274 => (x"78",x"c2",x"48",x"d0"),
   275 => (x"e4",x"f3",x"48",x"73"),
   276 => (x"5b",x"5e",x"0e",x"87"),
   277 => (x"c0",x"0e",x"5d",x"5c"),
   278 => (x"f0",x"ff",x"c0",x"1e"),
   279 => (x"f3",x"49",x"c9",x"c1"),
   280 => (x"1e",x"d2",x"87",x"d7"),
   281 => (x"49",x"f0",x"dc",x"c2"),
   282 => (x"c8",x"87",x"fd",x"fc"),
   283 => (x"c1",x"4c",x"c0",x"86"),
   284 => (x"ac",x"b7",x"d2",x"84"),
   285 => (x"c2",x"87",x"f8",x"04"),
   286 => (x"bf",x"97",x"f0",x"dc"),
   287 => (x"99",x"c0",x"c3",x"49"),
   288 => (x"05",x"a9",x"c0",x"c1"),
   289 => (x"c2",x"87",x"e7",x"c0"),
   290 => (x"bf",x"97",x"f7",x"dc"),
   291 => (x"c2",x"31",x"d0",x"49"),
   292 => (x"bf",x"97",x"f8",x"dc"),
   293 => (x"72",x"32",x"c8",x"4a"),
   294 => (x"f9",x"dc",x"c2",x"b1"),
   295 => (x"b1",x"4a",x"bf",x"97"),
   296 => (x"ff",x"cf",x"4c",x"71"),
   297 => (x"c1",x"9c",x"ff",x"ff"),
   298 => (x"c1",x"34",x"ca",x"84"),
   299 => (x"dc",x"c2",x"87",x"e7"),
   300 => (x"49",x"bf",x"97",x"f9"),
   301 => (x"99",x"c6",x"31",x"c1"),
   302 => (x"97",x"fa",x"dc",x"c2"),
   303 => (x"b7",x"c7",x"4a",x"bf"),
   304 => (x"c2",x"b1",x"72",x"2a"),
   305 => (x"bf",x"97",x"f5",x"dc"),
   306 => (x"9d",x"cf",x"4d",x"4a"),
   307 => (x"97",x"f6",x"dc",x"c2"),
   308 => (x"9a",x"c3",x"4a",x"bf"),
   309 => (x"dc",x"c2",x"32",x"ca"),
   310 => (x"4b",x"bf",x"97",x"f7"),
   311 => (x"b2",x"73",x"33",x"c2"),
   312 => (x"97",x"f8",x"dc",x"c2"),
   313 => (x"c0",x"c3",x"4b",x"bf"),
   314 => (x"2b",x"b7",x"c6",x"9b"),
   315 => (x"81",x"c2",x"b2",x"73"),
   316 => (x"30",x"71",x"48",x"c1"),
   317 => (x"48",x"c1",x"49",x"70"),
   318 => (x"4d",x"70",x"30",x"75"),
   319 => (x"84",x"c1",x"4c",x"72"),
   320 => (x"c0",x"c8",x"94",x"71"),
   321 => (x"cc",x"06",x"ad",x"b7"),
   322 => (x"b7",x"34",x"c1",x"87"),
   323 => (x"b7",x"c0",x"c8",x"2d"),
   324 => (x"f4",x"ff",x"01",x"ad"),
   325 => (x"f0",x"48",x"74",x"87"),
   326 => (x"5e",x"0e",x"87",x"d7"),
   327 => (x"0e",x"5d",x"5c",x"5b"),
   328 => (x"e5",x"c2",x"86",x"f8"),
   329 => (x"78",x"c0",x"48",x"d6"),
   330 => (x"1e",x"ce",x"dd",x"c2"),
   331 => (x"de",x"fb",x"49",x"c0"),
   332 => (x"70",x"86",x"c4",x"87"),
   333 => (x"87",x"c5",x"05",x"98"),
   334 => (x"c0",x"c9",x"48",x"c0"),
   335 => (x"c1",x"4d",x"c0",x"87"),
   336 => (x"dd",x"f2",x"c0",x"7e"),
   337 => (x"de",x"c2",x"49",x"bf"),
   338 => (x"c8",x"71",x"4a",x"c4"),
   339 => (x"87",x"d9",x"ec",x"4b"),
   340 => (x"c2",x"05",x"98",x"70"),
   341 => (x"c0",x"7e",x"c0",x"87"),
   342 => (x"49",x"bf",x"d9",x"f2"),
   343 => (x"4a",x"e0",x"de",x"c2"),
   344 => (x"ec",x"4b",x"c8",x"71"),
   345 => (x"98",x"70",x"87",x"c3"),
   346 => (x"c0",x"87",x"c2",x"05"),
   347 => (x"c0",x"02",x"6e",x"7e"),
   348 => (x"e4",x"c2",x"87",x"fd"),
   349 => (x"c2",x"4d",x"bf",x"d4"),
   350 => (x"bf",x"9f",x"cc",x"e5"),
   351 => (x"d6",x"c5",x"48",x"7e"),
   352 => (x"c7",x"05",x"a8",x"ea"),
   353 => (x"d4",x"e4",x"c2",x"87"),
   354 => (x"87",x"ce",x"4d",x"bf"),
   355 => (x"e9",x"ca",x"48",x"6e"),
   356 => (x"c5",x"02",x"a8",x"d5"),
   357 => (x"c7",x"48",x"c0",x"87"),
   358 => (x"dd",x"c2",x"87",x"e3"),
   359 => (x"49",x"75",x"1e",x"ce"),
   360 => (x"c4",x"87",x"ec",x"f9"),
   361 => (x"05",x"98",x"70",x"86"),
   362 => (x"48",x"c0",x"87",x"c5"),
   363 => (x"c0",x"87",x"ce",x"c7"),
   364 => (x"49",x"bf",x"d9",x"f2"),
   365 => (x"4a",x"e0",x"de",x"c2"),
   366 => (x"ea",x"4b",x"c8",x"71"),
   367 => (x"98",x"70",x"87",x"eb"),
   368 => (x"c2",x"87",x"c8",x"05"),
   369 => (x"c1",x"48",x"d6",x"e5"),
   370 => (x"c0",x"87",x"da",x"78"),
   371 => (x"49",x"bf",x"dd",x"f2"),
   372 => (x"4a",x"c4",x"de",x"c2"),
   373 => (x"ea",x"4b",x"c8",x"71"),
   374 => (x"98",x"70",x"87",x"cf"),
   375 => (x"87",x"c5",x"c0",x"02"),
   376 => (x"d8",x"c6",x"48",x"c0"),
   377 => (x"cc",x"e5",x"c2",x"87"),
   378 => (x"c1",x"49",x"bf",x"97"),
   379 => (x"c0",x"05",x"a9",x"d5"),
   380 => (x"e5",x"c2",x"87",x"cd"),
   381 => (x"49",x"bf",x"97",x"cd"),
   382 => (x"02",x"a9",x"ea",x"c2"),
   383 => (x"c0",x"87",x"c5",x"c0"),
   384 => (x"87",x"f9",x"c5",x"48"),
   385 => (x"97",x"ce",x"dd",x"c2"),
   386 => (x"c3",x"48",x"7e",x"bf"),
   387 => (x"c0",x"02",x"a8",x"e9"),
   388 => (x"48",x"6e",x"87",x"ce"),
   389 => (x"02",x"a8",x"eb",x"c3"),
   390 => (x"c0",x"87",x"c5",x"c0"),
   391 => (x"87",x"dd",x"c5",x"48"),
   392 => (x"97",x"d9",x"dd",x"c2"),
   393 => (x"05",x"99",x"49",x"bf"),
   394 => (x"c2",x"87",x"cc",x"c0"),
   395 => (x"bf",x"97",x"da",x"dd"),
   396 => (x"02",x"a9",x"c2",x"49"),
   397 => (x"c0",x"87",x"c5",x"c0"),
   398 => (x"87",x"c1",x"c5",x"48"),
   399 => (x"97",x"db",x"dd",x"c2"),
   400 => (x"e5",x"c2",x"48",x"bf"),
   401 => (x"4c",x"70",x"58",x"d2"),
   402 => (x"c2",x"88",x"c1",x"48"),
   403 => (x"c2",x"58",x"d6",x"e5"),
   404 => (x"bf",x"97",x"dc",x"dd"),
   405 => (x"c2",x"81",x"75",x"49"),
   406 => (x"bf",x"97",x"dd",x"dd"),
   407 => (x"72",x"32",x"c8",x"4a"),
   408 => (x"e9",x"c2",x"7e",x"a1"),
   409 => (x"78",x"6e",x"48",x"e3"),
   410 => (x"97",x"de",x"dd",x"c2"),
   411 => (x"a6",x"c8",x"48",x"bf"),
   412 => (x"d6",x"e5",x"c2",x"58"),
   413 => (x"cf",x"c2",x"02",x"bf"),
   414 => (x"d9",x"f2",x"c0",x"87"),
   415 => (x"de",x"c2",x"49",x"bf"),
   416 => (x"c8",x"71",x"4a",x"e0"),
   417 => (x"87",x"e1",x"e7",x"4b"),
   418 => (x"c0",x"02",x"98",x"70"),
   419 => (x"48",x"c0",x"87",x"c5"),
   420 => (x"c2",x"87",x"ea",x"c3"),
   421 => (x"4c",x"bf",x"ce",x"e5"),
   422 => (x"5c",x"f7",x"e9",x"c2"),
   423 => (x"97",x"f3",x"dd",x"c2"),
   424 => (x"31",x"c8",x"49",x"bf"),
   425 => (x"97",x"f2",x"dd",x"c2"),
   426 => (x"49",x"a1",x"4a",x"bf"),
   427 => (x"97",x"f4",x"dd",x"c2"),
   428 => (x"32",x"d0",x"4a",x"bf"),
   429 => (x"c2",x"49",x"a1",x"72"),
   430 => (x"bf",x"97",x"f5",x"dd"),
   431 => (x"72",x"32",x"d8",x"4a"),
   432 => (x"66",x"c4",x"49",x"a1"),
   433 => (x"e3",x"e9",x"c2",x"91"),
   434 => (x"e9",x"c2",x"81",x"bf"),
   435 => (x"dd",x"c2",x"59",x"eb"),
   436 => (x"4a",x"bf",x"97",x"fb"),
   437 => (x"dd",x"c2",x"32",x"c8"),
   438 => (x"4b",x"bf",x"97",x"fa"),
   439 => (x"dd",x"c2",x"4a",x"a2"),
   440 => (x"4b",x"bf",x"97",x"fc"),
   441 => (x"a2",x"73",x"33",x"d0"),
   442 => (x"fd",x"dd",x"c2",x"4a"),
   443 => (x"cf",x"4b",x"bf",x"97"),
   444 => (x"73",x"33",x"d8",x"9b"),
   445 => (x"e9",x"c2",x"4a",x"a2"),
   446 => (x"8a",x"c2",x"5a",x"ef"),
   447 => (x"e9",x"c2",x"92",x"74"),
   448 => (x"a1",x"72",x"48",x"ef"),
   449 => (x"87",x"c1",x"c1",x"78"),
   450 => (x"97",x"e0",x"dd",x"c2"),
   451 => (x"31",x"c8",x"49",x"bf"),
   452 => (x"97",x"df",x"dd",x"c2"),
   453 => (x"49",x"a1",x"4a",x"bf"),
   454 => (x"ff",x"c7",x"31",x"c5"),
   455 => (x"c2",x"29",x"c9",x"81"),
   456 => (x"c2",x"59",x"f7",x"e9"),
   457 => (x"bf",x"97",x"e5",x"dd"),
   458 => (x"c2",x"32",x"c8",x"4a"),
   459 => (x"bf",x"97",x"e4",x"dd"),
   460 => (x"c4",x"4a",x"a2",x"4b"),
   461 => (x"82",x"6e",x"92",x"66"),
   462 => (x"5a",x"f3",x"e9",x"c2"),
   463 => (x"48",x"eb",x"e9",x"c2"),
   464 => (x"e9",x"c2",x"78",x"c0"),
   465 => (x"a1",x"72",x"48",x"e7"),
   466 => (x"f7",x"e9",x"c2",x"78"),
   467 => (x"eb",x"e9",x"c2",x"48"),
   468 => (x"e9",x"c2",x"78",x"bf"),
   469 => (x"e9",x"c2",x"48",x"fb"),
   470 => (x"c2",x"78",x"bf",x"ef"),
   471 => (x"02",x"bf",x"d6",x"e5"),
   472 => (x"74",x"87",x"c9",x"c0"),
   473 => (x"70",x"30",x"c4",x"48"),
   474 => (x"87",x"c9",x"c0",x"7e"),
   475 => (x"bf",x"f3",x"e9",x"c2"),
   476 => (x"70",x"30",x"c4",x"48"),
   477 => (x"da",x"e5",x"c2",x"7e"),
   478 => (x"c1",x"78",x"6e",x"48"),
   479 => (x"26",x"8e",x"f8",x"48"),
   480 => (x"26",x"4c",x"26",x"4d"),
   481 => (x"0e",x"4f",x"26",x"4b"),
   482 => (x"5d",x"5c",x"5b",x"5e"),
   483 => (x"c2",x"4a",x"71",x"0e"),
   484 => (x"02",x"bf",x"d6",x"e5"),
   485 => (x"4b",x"72",x"87",x"cb"),
   486 => (x"4d",x"72",x"2b",x"c7"),
   487 => (x"c9",x"9d",x"ff",x"c1"),
   488 => (x"c8",x"4b",x"72",x"87"),
   489 => (x"c3",x"4d",x"72",x"2b"),
   490 => (x"e9",x"c2",x"9d",x"ff"),
   491 => (x"c0",x"83",x"bf",x"e3"),
   492 => (x"ab",x"bf",x"d5",x"f2"),
   493 => (x"c0",x"87",x"d9",x"02"),
   494 => (x"c2",x"5b",x"d9",x"f2"),
   495 => (x"73",x"1e",x"ce",x"dd"),
   496 => (x"87",x"cb",x"f1",x"49"),
   497 => (x"98",x"70",x"86",x"c4"),
   498 => (x"c0",x"87",x"c5",x"05"),
   499 => (x"87",x"e6",x"c0",x"48"),
   500 => (x"bf",x"d6",x"e5",x"c2"),
   501 => (x"75",x"87",x"d2",x"02"),
   502 => (x"c2",x"91",x"c4",x"49"),
   503 => (x"69",x"81",x"ce",x"dd"),
   504 => (x"ff",x"ff",x"cf",x"4c"),
   505 => (x"cb",x"9c",x"ff",x"ff"),
   506 => (x"c2",x"49",x"75",x"87"),
   507 => (x"ce",x"dd",x"c2",x"91"),
   508 => (x"4c",x"69",x"9f",x"81"),
   509 => (x"c6",x"fe",x"48",x"74"),
   510 => (x"5b",x"5e",x"0e",x"87"),
   511 => (x"f8",x"0e",x"5d",x"5c"),
   512 => (x"9c",x"4c",x"71",x"86"),
   513 => (x"c0",x"87",x"c5",x"05"),
   514 => (x"87",x"c0",x"c3",x"48"),
   515 => (x"48",x"7e",x"a4",x"c8"),
   516 => (x"66",x"d8",x"78",x"c0"),
   517 => (x"d8",x"87",x"c7",x"02"),
   518 => (x"05",x"bf",x"97",x"66"),
   519 => (x"48",x"c0",x"87",x"c5"),
   520 => (x"c0",x"87",x"e9",x"c2"),
   521 => (x"49",x"49",x"c1",x"1e"),
   522 => (x"c4",x"87",x"d3",x"ca"),
   523 => (x"9d",x"4d",x"70",x"86"),
   524 => (x"87",x"c2",x"c1",x"02"),
   525 => (x"4a",x"de",x"e5",x"c2"),
   526 => (x"e0",x"49",x"66",x"d8"),
   527 => (x"98",x"70",x"87",x"d0"),
   528 => (x"87",x"f2",x"c0",x"02"),
   529 => (x"66",x"d8",x"4a",x"75"),
   530 => (x"e0",x"4b",x"cb",x"49"),
   531 => (x"98",x"70",x"87",x"f5"),
   532 => (x"87",x"e2",x"c0",x"02"),
   533 => (x"9d",x"75",x"1e",x"c0"),
   534 => (x"c8",x"87",x"c7",x"02"),
   535 => (x"78",x"c0",x"48",x"a6"),
   536 => (x"a6",x"c8",x"87",x"c5"),
   537 => (x"c8",x"78",x"c1",x"48"),
   538 => (x"d1",x"c9",x"49",x"66"),
   539 => (x"70",x"86",x"c4",x"87"),
   540 => (x"fe",x"05",x"9d",x"4d"),
   541 => (x"9d",x"75",x"87",x"fe"),
   542 => (x"87",x"ce",x"c1",x"02"),
   543 => (x"6e",x"49",x"a5",x"dc"),
   544 => (x"da",x"78",x"69",x"48"),
   545 => (x"a6",x"c4",x"49",x"a5"),
   546 => (x"78",x"a4",x"c4",x"48"),
   547 => (x"c4",x"48",x"69",x"9f"),
   548 => (x"c2",x"78",x"08",x"66"),
   549 => (x"02",x"bf",x"d6",x"e5"),
   550 => (x"a5",x"d4",x"87",x"d2"),
   551 => (x"49",x"69",x"9f",x"49"),
   552 => (x"99",x"ff",x"ff",x"c0"),
   553 => (x"30",x"d0",x"48",x"71"),
   554 => (x"87",x"c2",x"7e",x"70"),
   555 => (x"48",x"6e",x"7e",x"c0"),
   556 => (x"80",x"bf",x"66",x"c4"),
   557 => (x"78",x"08",x"66",x"c4"),
   558 => (x"a4",x"cc",x"7c",x"c0"),
   559 => (x"bf",x"66",x"c4",x"49"),
   560 => (x"49",x"a4",x"d0",x"79"),
   561 => (x"48",x"c1",x"79",x"c0"),
   562 => (x"48",x"c0",x"87",x"c2"),
   563 => (x"ee",x"fa",x"8e",x"f8"),
   564 => (x"5b",x"5e",x"0e",x"87"),
   565 => (x"4c",x"71",x"0e",x"5c"),
   566 => (x"cb",x"c1",x"02",x"9c"),
   567 => (x"49",x"a4",x"c8",x"87"),
   568 => (x"c3",x"c1",x"02",x"69"),
   569 => (x"cc",x"49",x"6c",x"87"),
   570 => (x"80",x"71",x"48",x"66"),
   571 => (x"70",x"58",x"a6",x"d0"),
   572 => (x"d2",x"e5",x"c2",x"b9"),
   573 => (x"ba",x"ff",x"4a",x"bf"),
   574 => (x"99",x"71",x"99",x"72"),
   575 => (x"87",x"e5",x"c0",x"02"),
   576 => (x"6b",x"4b",x"a4",x"c4"),
   577 => (x"87",x"ff",x"f9",x"49"),
   578 => (x"e5",x"c2",x"7b",x"70"),
   579 => (x"6c",x"49",x"bf",x"ce"),
   580 => (x"cc",x"7c",x"71",x"81"),
   581 => (x"e5",x"c2",x"b9",x"66"),
   582 => (x"ff",x"4a",x"bf",x"d2"),
   583 => (x"71",x"99",x"72",x"ba"),
   584 => (x"db",x"ff",x"05",x"99"),
   585 => (x"7c",x"66",x"cc",x"87"),
   586 => (x"1e",x"87",x"d6",x"f9"),
   587 => (x"4b",x"71",x"1e",x"73"),
   588 => (x"87",x"c7",x"02",x"9b"),
   589 => (x"69",x"49",x"a3",x"c8"),
   590 => (x"c0",x"87",x"c5",x"05"),
   591 => (x"87",x"f6",x"c0",x"48"),
   592 => (x"bf",x"e7",x"e9",x"c2"),
   593 => (x"4a",x"a3",x"c4",x"49"),
   594 => (x"8a",x"c2",x"4a",x"6a"),
   595 => (x"bf",x"ce",x"e5",x"c2"),
   596 => (x"49",x"a1",x"72",x"92"),
   597 => (x"bf",x"d2",x"e5",x"c2"),
   598 => (x"72",x"9a",x"6b",x"4a"),
   599 => (x"f2",x"c0",x"49",x"a1"),
   600 => (x"66",x"c8",x"59",x"d9"),
   601 => (x"e6",x"ea",x"71",x"1e"),
   602 => (x"70",x"86",x"c4",x"87"),
   603 => (x"87",x"c4",x"05",x"98"),
   604 => (x"87",x"c2",x"48",x"c0"),
   605 => (x"ca",x"f8",x"48",x"c1"),
   606 => (x"1e",x"73",x"1e",x"87"),
   607 => (x"02",x"9b",x"4b",x"71"),
   608 => (x"a3",x"c8",x"87",x"c7"),
   609 => (x"c5",x"05",x"69",x"49"),
   610 => (x"c0",x"48",x"c0",x"87"),
   611 => (x"e9",x"c2",x"87",x"f6"),
   612 => (x"c4",x"49",x"bf",x"e7"),
   613 => (x"4a",x"6a",x"4a",x"a3"),
   614 => (x"e5",x"c2",x"8a",x"c2"),
   615 => (x"72",x"92",x"bf",x"ce"),
   616 => (x"e5",x"c2",x"49",x"a1"),
   617 => (x"6b",x"4a",x"bf",x"d2"),
   618 => (x"49",x"a1",x"72",x"9a"),
   619 => (x"59",x"d9",x"f2",x"c0"),
   620 => (x"71",x"1e",x"66",x"c8"),
   621 => (x"c4",x"87",x"d1",x"e6"),
   622 => (x"05",x"98",x"70",x"86"),
   623 => (x"48",x"c0",x"87",x"c4"),
   624 => (x"48",x"c1",x"87",x"c2"),
   625 => (x"0e",x"87",x"fc",x"f6"),
   626 => (x"5d",x"5c",x"5b",x"5e"),
   627 => (x"4b",x"71",x"1e",x"0e"),
   628 => (x"73",x"4d",x"66",x"d4"),
   629 => (x"cc",x"c1",x"02",x"9b"),
   630 => (x"49",x"a3",x"c8",x"87"),
   631 => (x"c4",x"c1",x"02",x"69"),
   632 => (x"4c",x"a3",x"d0",x"87"),
   633 => (x"bf",x"d2",x"e5",x"c2"),
   634 => (x"6c",x"b9",x"ff",x"49"),
   635 => (x"d4",x"7e",x"99",x"4a"),
   636 => (x"cd",x"06",x"a9",x"66"),
   637 => (x"7c",x"7b",x"c0",x"87"),
   638 => (x"c4",x"4a",x"a3",x"cc"),
   639 => (x"79",x"6a",x"49",x"a3"),
   640 => (x"49",x"72",x"87",x"ca"),
   641 => (x"d4",x"99",x"c0",x"f8"),
   642 => (x"8d",x"71",x"4d",x"66"),
   643 => (x"29",x"c9",x"49",x"75"),
   644 => (x"49",x"73",x"1e",x"71"),
   645 => (x"c2",x"87",x"fa",x"fa"),
   646 => (x"73",x"1e",x"ce",x"dd"),
   647 => (x"87",x"cb",x"fc",x"49"),
   648 => (x"66",x"d4",x"86",x"c8"),
   649 => (x"d6",x"f5",x"26",x"7c"),
   650 => (x"1e",x"73",x"1e",x"87"),
   651 => (x"02",x"9b",x"4b",x"71"),
   652 => (x"c2",x"87",x"e4",x"c0"),
   653 => (x"73",x"5b",x"fb",x"e9"),
   654 => (x"c2",x"8a",x"c2",x"4a"),
   655 => (x"49",x"bf",x"ce",x"e5"),
   656 => (x"e7",x"e9",x"c2",x"92"),
   657 => (x"80",x"72",x"48",x"bf"),
   658 => (x"58",x"ff",x"e9",x"c2"),
   659 => (x"30",x"c4",x"48",x"71"),
   660 => (x"58",x"de",x"e5",x"c2"),
   661 => (x"c2",x"87",x"ed",x"c0"),
   662 => (x"c2",x"48",x"f7",x"e9"),
   663 => (x"78",x"bf",x"eb",x"e9"),
   664 => (x"48",x"fb",x"e9",x"c2"),
   665 => (x"bf",x"ef",x"e9",x"c2"),
   666 => (x"d6",x"e5",x"c2",x"78"),
   667 => (x"87",x"c9",x"02",x"bf"),
   668 => (x"bf",x"ce",x"e5",x"c2"),
   669 => (x"c7",x"31",x"c4",x"49"),
   670 => (x"f3",x"e9",x"c2",x"87"),
   671 => (x"31",x"c4",x"49",x"bf"),
   672 => (x"59",x"de",x"e5",x"c2"),
   673 => (x"0e",x"87",x"fc",x"f3"),
   674 => (x"0e",x"5c",x"5b",x"5e"),
   675 => (x"4b",x"c0",x"4a",x"71"),
   676 => (x"c0",x"02",x"9a",x"72"),
   677 => (x"a2",x"da",x"87",x"e0"),
   678 => (x"4b",x"69",x"9f",x"49"),
   679 => (x"bf",x"d6",x"e5",x"c2"),
   680 => (x"d4",x"87",x"cf",x"02"),
   681 => (x"69",x"9f",x"49",x"a2"),
   682 => (x"ff",x"c0",x"4c",x"49"),
   683 => (x"34",x"d0",x"9c",x"ff"),
   684 => (x"4c",x"c0",x"87",x"c2"),
   685 => (x"49",x"73",x"b3",x"74"),
   686 => (x"f3",x"87",x"ee",x"fd"),
   687 => (x"5e",x"0e",x"87",x"c3"),
   688 => (x"0e",x"5d",x"5c",x"5b"),
   689 => (x"4a",x"71",x"86",x"f4"),
   690 => (x"9a",x"72",x"7e",x"c0"),
   691 => (x"c2",x"87",x"d8",x"02"),
   692 => (x"c0",x"48",x"ca",x"dd"),
   693 => (x"c2",x"dd",x"c2",x"78"),
   694 => (x"fb",x"e9",x"c2",x"48"),
   695 => (x"dd",x"c2",x"78",x"bf"),
   696 => (x"e9",x"c2",x"48",x"c6"),
   697 => (x"c2",x"78",x"bf",x"f7"),
   698 => (x"c0",x"48",x"eb",x"e5"),
   699 => (x"da",x"e5",x"c2",x"50"),
   700 => (x"dd",x"c2",x"49",x"bf"),
   701 => (x"71",x"4a",x"bf",x"ca"),
   702 => (x"c9",x"c4",x"03",x"aa"),
   703 => (x"cf",x"49",x"72",x"87"),
   704 => (x"e9",x"c0",x"05",x"99"),
   705 => (x"d5",x"f2",x"c0",x"87"),
   706 => (x"c2",x"dd",x"c2",x"48"),
   707 => (x"dd",x"c2",x"78",x"bf"),
   708 => (x"dd",x"c2",x"1e",x"ce"),
   709 => (x"c2",x"49",x"bf",x"c2"),
   710 => (x"c1",x"48",x"c2",x"dd"),
   711 => (x"e3",x"71",x"78",x"a1"),
   712 => (x"86",x"c4",x"87",x"ed"),
   713 => (x"48",x"d1",x"f2",x"c0"),
   714 => (x"78",x"ce",x"dd",x"c2"),
   715 => (x"f2",x"c0",x"87",x"cc"),
   716 => (x"c0",x"48",x"bf",x"d1"),
   717 => (x"f2",x"c0",x"80",x"e0"),
   718 => (x"dd",x"c2",x"58",x"d5"),
   719 => (x"c1",x"48",x"bf",x"ca"),
   720 => (x"ce",x"dd",x"c2",x"80"),
   721 => (x"0c",x"91",x"27",x"58"),
   722 => (x"97",x"bf",x"00",x"00"),
   723 => (x"02",x"9d",x"4d",x"bf"),
   724 => (x"c3",x"87",x"e3",x"c2"),
   725 => (x"c2",x"02",x"ad",x"e5"),
   726 => (x"f2",x"c0",x"87",x"dc"),
   727 => (x"cb",x"4b",x"bf",x"d1"),
   728 => (x"4c",x"11",x"49",x"a3"),
   729 => (x"c1",x"05",x"ac",x"cf"),
   730 => (x"49",x"75",x"87",x"d2"),
   731 => (x"89",x"c1",x"99",x"df"),
   732 => (x"e5",x"c2",x"91",x"cd"),
   733 => (x"a3",x"c1",x"81",x"de"),
   734 => (x"c3",x"51",x"12",x"4a"),
   735 => (x"51",x"12",x"4a",x"a3"),
   736 => (x"12",x"4a",x"a3",x"c5"),
   737 => (x"4a",x"a3",x"c7",x"51"),
   738 => (x"a3",x"c9",x"51",x"12"),
   739 => (x"ce",x"51",x"12",x"4a"),
   740 => (x"51",x"12",x"4a",x"a3"),
   741 => (x"12",x"4a",x"a3",x"d0"),
   742 => (x"4a",x"a3",x"d2",x"51"),
   743 => (x"a3",x"d4",x"51",x"12"),
   744 => (x"d6",x"51",x"12",x"4a"),
   745 => (x"51",x"12",x"4a",x"a3"),
   746 => (x"12",x"4a",x"a3",x"d8"),
   747 => (x"4a",x"a3",x"dc",x"51"),
   748 => (x"a3",x"de",x"51",x"12"),
   749 => (x"c1",x"51",x"12",x"4a"),
   750 => (x"87",x"fa",x"c0",x"7e"),
   751 => (x"99",x"c8",x"49",x"74"),
   752 => (x"87",x"eb",x"c0",x"05"),
   753 => (x"99",x"d0",x"49",x"74"),
   754 => (x"dc",x"87",x"d1",x"05"),
   755 => (x"cb",x"c0",x"02",x"66"),
   756 => (x"dc",x"49",x"73",x"87"),
   757 => (x"98",x"70",x"0f",x"66"),
   758 => (x"87",x"d3",x"c0",x"02"),
   759 => (x"c6",x"c0",x"05",x"6e"),
   760 => (x"de",x"e5",x"c2",x"87"),
   761 => (x"c0",x"50",x"c0",x"48"),
   762 => (x"48",x"bf",x"d1",x"f2"),
   763 => (x"c2",x"87",x"dd",x"c2"),
   764 => (x"c0",x"48",x"eb",x"e5"),
   765 => (x"e5",x"c2",x"7e",x"50"),
   766 => (x"c2",x"49",x"bf",x"da"),
   767 => (x"4a",x"bf",x"ca",x"dd"),
   768 => (x"fb",x"04",x"aa",x"71"),
   769 => (x"e9",x"c2",x"87",x"f7"),
   770 => (x"c0",x"05",x"bf",x"fb"),
   771 => (x"e5",x"c2",x"87",x"c8"),
   772 => (x"c1",x"02",x"bf",x"d6"),
   773 => (x"dd",x"c2",x"87",x"f4"),
   774 => (x"ed",x"49",x"bf",x"c6"),
   775 => (x"dd",x"c2",x"87",x"e9"),
   776 => (x"a6",x"c4",x"58",x"ca"),
   777 => (x"c6",x"dd",x"c2",x"48"),
   778 => (x"e5",x"c2",x"78",x"bf"),
   779 => (x"c0",x"02",x"bf",x"d6"),
   780 => (x"66",x"c4",x"87",x"d8"),
   781 => (x"ff",x"ff",x"cf",x"49"),
   782 => (x"a9",x"99",x"f8",x"ff"),
   783 => (x"87",x"c5",x"c0",x"02"),
   784 => (x"e1",x"c0",x"4c",x"c0"),
   785 => (x"c0",x"4c",x"c1",x"87"),
   786 => (x"66",x"c4",x"87",x"dc"),
   787 => (x"f8",x"ff",x"cf",x"49"),
   788 => (x"c0",x"02",x"a9",x"99"),
   789 => (x"a6",x"c8",x"87",x"c8"),
   790 => (x"c0",x"78",x"c0",x"48"),
   791 => (x"a6",x"c8",x"87",x"c5"),
   792 => (x"c8",x"78",x"c1",x"48"),
   793 => (x"9c",x"74",x"4c",x"66"),
   794 => (x"87",x"de",x"c0",x"05"),
   795 => (x"c2",x"49",x"66",x"c4"),
   796 => (x"ce",x"e5",x"c2",x"89"),
   797 => (x"e9",x"c2",x"91",x"bf"),
   798 => (x"71",x"48",x"bf",x"e7"),
   799 => (x"c6",x"dd",x"c2",x"80"),
   800 => (x"ca",x"dd",x"c2",x"58"),
   801 => (x"f9",x"78",x"c0",x"48"),
   802 => (x"48",x"c0",x"87",x"e3"),
   803 => (x"ee",x"eb",x"8e",x"f4"),
   804 => (x"00",x"00",x"00",x"87"),
   805 => (x"ff",x"ff",x"ff",x"00"),
   806 => (x"00",x"0c",x"a1",x"ff"),
   807 => (x"00",x"0c",x"aa",x"00"),
   808 => (x"54",x"41",x"46",x"00"),
   809 => (x"20",x"20",x"32",x"33"),
   810 => (x"41",x"46",x"00",x"20"),
   811 => (x"20",x"36",x"31",x"54"),
   812 => (x"1e",x"00",x"20",x"20"),
   813 => (x"c3",x"48",x"d4",x"ff"),
   814 => (x"48",x"68",x"78",x"ff"),
   815 => (x"ff",x"1e",x"4f",x"26"),
   816 => (x"ff",x"c3",x"48",x"d4"),
   817 => (x"48",x"d0",x"ff",x"78"),
   818 => (x"ff",x"78",x"e1",x"c0"),
   819 => (x"78",x"d4",x"48",x"d4"),
   820 => (x"48",x"ff",x"e9",x"c2"),
   821 => (x"50",x"bf",x"d4",x"ff"),
   822 => (x"ff",x"1e",x"4f",x"26"),
   823 => (x"e0",x"c0",x"48",x"d0"),
   824 => (x"1e",x"4f",x"26",x"78"),
   825 => (x"70",x"87",x"cc",x"ff"),
   826 => (x"c6",x"02",x"99",x"49"),
   827 => (x"a9",x"fb",x"c0",x"87"),
   828 => (x"71",x"87",x"f1",x"05"),
   829 => (x"0e",x"4f",x"26",x"48"),
   830 => (x"0e",x"5c",x"5b",x"5e"),
   831 => (x"4c",x"c0",x"4b",x"71"),
   832 => (x"70",x"87",x"f0",x"fe"),
   833 => (x"c0",x"02",x"99",x"49"),
   834 => (x"ec",x"c0",x"87",x"f9"),
   835 => (x"f2",x"c0",x"02",x"a9"),
   836 => (x"a9",x"fb",x"c0",x"87"),
   837 => (x"87",x"eb",x"c0",x"02"),
   838 => (x"ac",x"b7",x"66",x"cc"),
   839 => (x"d0",x"87",x"c7",x"03"),
   840 => (x"87",x"c2",x"02",x"66"),
   841 => (x"99",x"71",x"53",x"71"),
   842 => (x"c1",x"87",x"c2",x"02"),
   843 => (x"87",x"c3",x"fe",x"84"),
   844 => (x"02",x"99",x"49",x"70"),
   845 => (x"ec",x"c0",x"87",x"cd"),
   846 => (x"87",x"c7",x"02",x"a9"),
   847 => (x"05",x"a9",x"fb",x"c0"),
   848 => (x"d0",x"87",x"d5",x"ff"),
   849 => (x"87",x"c3",x"02",x"66"),
   850 => (x"c0",x"7b",x"97",x"c0"),
   851 => (x"c4",x"05",x"a9",x"ec"),
   852 => (x"c5",x"4a",x"74",x"87"),
   853 => (x"c0",x"4a",x"74",x"87"),
   854 => (x"48",x"72",x"8a",x"0a"),
   855 => (x"4d",x"26",x"87",x"c2"),
   856 => (x"4b",x"26",x"4c",x"26"),
   857 => (x"fd",x"1e",x"4f",x"26"),
   858 => (x"49",x"70",x"87",x"c9"),
   859 => (x"aa",x"f0",x"c0",x"4a"),
   860 => (x"c0",x"87",x"c9",x"04"),
   861 => (x"c3",x"01",x"aa",x"f9"),
   862 => (x"8a",x"f0",x"c0",x"87"),
   863 => (x"04",x"aa",x"c1",x"c1"),
   864 => (x"da",x"c1",x"87",x"c9"),
   865 => (x"87",x"c3",x"01",x"aa"),
   866 => (x"72",x"8a",x"f7",x"c0"),
   867 => (x"0e",x"4f",x"26",x"48"),
   868 => (x"5d",x"5c",x"5b",x"5e"),
   869 => (x"71",x"86",x"f8",x"0e"),
   870 => (x"fc",x"4d",x"c0",x"4c"),
   871 => (x"4b",x"c0",x"87",x"e0"),
   872 => (x"97",x"ee",x"f8",x"c0"),
   873 => (x"a9",x"c0",x"49",x"bf"),
   874 => (x"fc",x"87",x"cf",x"04"),
   875 => (x"83",x"c1",x"87",x"f5"),
   876 => (x"97",x"ee",x"f8",x"c0"),
   877 => (x"06",x"ab",x"49",x"bf"),
   878 => (x"f8",x"c0",x"87",x"f1"),
   879 => (x"02",x"bf",x"97",x"ee"),
   880 => (x"ee",x"fb",x"87",x"cf"),
   881 => (x"99",x"49",x"70",x"87"),
   882 => (x"c0",x"87",x"c6",x"02"),
   883 => (x"f1",x"05",x"a9",x"ec"),
   884 => (x"fb",x"4b",x"c0",x"87"),
   885 => (x"7e",x"70",x"87",x"dd"),
   886 => (x"c8",x"87",x"d8",x"fb"),
   887 => (x"d2",x"fb",x"58",x"a6"),
   888 => (x"c1",x"4a",x"70",x"87"),
   889 => (x"49",x"a4",x"c8",x"83"),
   890 => (x"6e",x"49",x"69",x"97"),
   891 => (x"87",x"da",x"05",x"a9"),
   892 => (x"97",x"49",x"a4",x"c9"),
   893 => (x"66",x"c4",x"49",x"69"),
   894 => (x"87",x"ce",x"05",x"a9"),
   895 => (x"97",x"49",x"a4",x"ca"),
   896 => (x"05",x"aa",x"49",x"69"),
   897 => (x"4d",x"c1",x"87",x"c4"),
   898 => (x"48",x"6e",x"87",x"d4"),
   899 => (x"02",x"a8",x"ec",x"c0"),
   900 => (x"48",x"6e",x"87",x"c8"),
   901 => (x"05",x"a8",x"fb",x"c0"),
   902 => (x"4b",x"c0",x"87",x"c4"),
   903 => (x"9d",x"75",x"4d",x"c1"),
   904 => (x"87",x"ef",x"fe",x"02"),
   905 => (x"73",x"87",x"f3",x"fa"),
   906 => (x"fc",x"8e",x"f8",x"48"),
   907 => (x"0e",x"00",x"87",x"f0"),
   908 => (x"5d",x"5c",x"5b",x"5e"),
   909 => (x"71",x"86",x"f8",x"0e"),
   910 => (x"4b",x"d4",x"ff",x"7e"),
   911 => (x"ea",x"c2",x"1e",x"6e"),
   912 => (x"f4",x"e6",x"49",x"c4"),
   913 => (x"70",x"86",x"c4",x"87"),
   914 => (x"ea",x"c4",x"02",x"98"),
   915 => (x"c2",x"e3",x"c1",x"87"),
   916 => (x"49",x"6e",x"4d",x"bf"),
   917 => (x"c8",x"87",x"f8",x"fc"),
   918 => (x"98",x"70",x"58",x"a6"),
   919 => (x"c4",x"87",x"c5",x"05"),
   920 => (x"78",x"c1",x"48",x"a6"),
   921 => (x"c5",x"48",x"d0",x"ff"),
   922 => (x"7b",x"d5",x"c1",x"78"),
   923 => (x"c1",x"49",x"66",x"c4"),
   924 => (x"c1",x"31",x"c6",x"89"),
   925 => (x"bf",x"97",x"c0",x"e3"),
   926 => (x"b0",x"71",x"48",x"4a"),
   927 => (x"d0",x"ff",x"7b",x"70"),
   928 => (x"c2",x"78",x"c4",x"48"),
   929 => (x"bf",x"97",x"ff",x"e9"),
   930 => (x"02",x"99",x"d0",x"49"),
   931 => (x"78",x"c5",x"87",x"d7"),
   932 => (x"c0",x"7b",x"d6",x"c1"),
   933 => (x"7b",x"ff",x"c3",x"4a"),
   934 => (x"e0",x"c0",x"82",x"c1"),
   935 => (x"87",x"f5",x"04",x"aa"),
   936 => (x"c4",x"48",x"d0",x"ff"),
   937 => (x"7b",x"ff",x"c3",x"78"),
   938 => (x"c5",x"48",x"d0",x"ff"),
   939 => (x"7b",x"d3",x"c1",x"78"),
   940 => (x"78",x"c4",x"7b",x"c1"),
   941 => (x"06",x"ad",x"b7",x"c0"),
   942 => (x"c2",x"87",x"eb",x"c2"),
   943 => (x"4c",x"bf",x"cc",x"ea"),
   944 => (x"c2",x"02",x"9c",x"8d"),
   945 => (x"dd",x"c2",x"87",x"c2"),
   946 => (x"a6",x"c4",x"7e",x"ce"),
   947 => (x"78",x"c0",x"c8",x"48"),
   948 => (x"ac",x"b7",x"c0",x"8c"),
   949 => (x"c8",x"87",x"c6",x"03"),
   950 => (x"c0",x"78",x"a4",x"c0"),
   951 => (x"ff",x"e9",x"c2",x"4c"),
   952 => (x"d0",x"49",x"bf",x"97"),
   953 => (x"87",x"d0",x"02",x"99"),
   954 => (x"ea",x"c2",x"1e",x"c0"),
   955 => (x"fa",x"e8",x"49",x"c4"),
   956 => (x"70",x"86",x"c4",x"87"),
   957 => (x"87",x"f5",x"c0",x"4a"),
   958 => (x"1e",x"ce",x"dd",x"c2"),
   959 => (x"49",x"c4",x"ea",x"c2"),
   960 => (x"c4",x"87",x"e8",x"e8"),
   961 => (x"ff",x"4a",x"70",x"86"),
   962 => (x"c5",x"c8",x"48",x"d0"),
   963 => (x"7b",x"d4",x"c1",x"78"),
   964 => (x"7b",x"bf",x"97",x"6e"),
   965 => (x"80",x"c1",x"48",x"6e"),
   966 => (x"66",x"c4",x"7e",x"70"),
   967 => (x"c8",x"88",x"c1",x"48"),
   968 => (x"98",x"70",x"58",x"a6"),
   969 => (x"87",x"e8",x"ff",x"05"),
   970 => (x"c4",x"48",x"d0",x"ff"),
   971 => (x"05",x"9a",x"72",x"78"),
   972 => (x"48",x"c0",x"87",x"c5"),
   973 => (x"c1",x"87",x"c2",x"c1"),
   974 => (x"c4",x"ea",x"c2",x"1e"),
   975 => (x"87",x"d1",x"e6",x"49"),
   976 => (x"9c",x"74",x"86",x"c4"),
   977 => (x"87",x"fe",x"fd",x"05"),
   978 => (x"06",x"ad",x"b7",x"c0"),
   979 => (x"ea",x"c2",x"87",x"d1"),
   980 => (x"78",x"c0",x"48",x"c4"),
   981 => (x"78",x"c0",x"80",x"d0"),
   982 => (x"ea",x"c2",x"80",x"f4"),
   983 => (x"c0",x"78",x"bf",x"d0"),
   984 => (x"fd",x"01",x"ad",x"b7"),
   985 => (x"d0",x"ff",x"87",x"d5"),
   986 => (x"c1",x"78",x"c5",x"48"),
   987 => (x"7b",x"c0",x"7b",x"d3"),
   988 => (x"48",x"c1",x"78",x"c4"),
   989 => (x"c0",x"87",x"c2",x"c0"),
   990 => (x"26",x"8e",x"f8",x"48"),
   991 => (x"26",x"4c",x"26",x"4d"),
   992 => (x"0e",x"4f",x"26",x"4b"),
   993 => (x"5d",x"5c",x"5b",x"5e"),
   994 => (x"4b",x"71",x"1e",x"0e"),
   995 => (x"ab",x"4d",x"4c",x"c0"),
   996 => (x"87",x"e8",x"c0",x"04"),
   997 => (x"1e",x"cf",x"f6",x"c0"),
   998 => (x"c4",x"02",x"9d",x"75"),
   999 => (x"c2",x"4a",x"c0",x"87"),
  1000 => (x"72",x"4a",x"c1",x"87"),
  1001 => (x"87",x"d6",x"ec",x"49"),
  1002 => (x"7e",x"70",x"86",x"c4"),
  1003 => (x"05",x"6e",x"84",x"c1"),
  1004 => (x"4c",x"73",x"87",x"c2"),
  1005 => (x"ac",x"73",x"85",x"c1"),
  1006 => (x"87",x"d8",x"ff",x"06"),
  1007 => (x"fe",x"26",x"48",x"6e"),
  1008 => (x"5e",x"0e",x"87",x"f9"),
  1009 => (x"71",x"0e",x"5c",x"5b"),
  1010 => (x"02",x"66",x"cc",x"4b"),
  1011 => (x"c0",x"4c",x"87",x"d8"),
  1012 => (x"d8",x"02",x"8c",x"f0"),
  1013 => (x"c1",x"4a",x"74",x"87"),
  1014 => (x"87",x"d1",x"02",x"8a"),
  1015 => (x"87",x"cd",x"02",x"8a"),
  1016 => (x"87",x"c9",x"02",x"8a"),
  1017 => (x"49",x"73",x"87",x"d9"),
  1018 => (x"d2",x"87",x"c4",x"f9"),
  1019 => (x"c0",x"1e",x"74",x"87"),
  1020 => (x"d4",x"d9",x"c1",x"49"),
  1021 => (x"73",x"1e",x"74",x"87"),
  1022 => (x"cc",x"d9",x"c1",x"49"),
  1023 => (x"fd",x"86",x"c8",x"87"),
  1024 => (x"5e",x"0e",x"87",x"fb"),
  1025 => (x"0e",x"5d",x"5c",x"5b"),
  1026 => (x"49",x"4c",x"71",x"1e"),
  1027 => (x"ea",x"c2",x"91",x"de"),
  1028 => (x"85",x"71",x"4d",x"ec"),
  1029 => (x"c1",x"02",x"6d",x"97"),
  1030 => (x"ea",x"c2",x"87",x"dc"),
  1031 => (x"74",x"49",x"bf",x"d8"),
  1032 => (x"de",x"fd",x"71",x"81"),
  1033 => (x"48",x"7e",x"70",x"87"),
  1034 => (x"f2",x"c0",x"02",x"98"),
  1035 => (x"e0",x"ea",x"c2",x"87"),
  1036 => (x"cb",x"4a",x"70",x"4b"),
  1037 => (x"ee",x"c1",x"ff",x"49"),
  1038 => (x"cb",x"4b",x"74",x"87"),
  1039 => (x"d4",x"e3",x"c1",x"93"),
  1040 => (x"c1",x"83",x"c4",x"83"),
  1041 => (x"74",x"7b",x"fa",x"c1"),
  1042 => (x"e4",x"c0",x"c1",x"49"),
  1043 => (x"c1",x"7b",x"75",x"87"),
  1044 => (x"bf",x"97",x"c1",x"e3"),
  1045 => (x"ea",x"c2",x"1e",x"49"),
  1046 => (x"e5",x"fd",x"49",x"e0"),
  1047 => (x"74",x"86",x"c4",x"87"),
  1048 => (x"cc",x"c0",x"c1",x"49"),
  1049 => (x"c1",x"49",x"c0",x"87"),
  1050 => (x"c2",x"87",x"eb",x"c1"),
  1051 => (x"c0",x"48",x"c0",x"ea"),
  1052 => (x"de",x"49",x"c1",x"78"),
  1053 => (x"fc",x"26",x"87",x"ca"),
  1054 => (x"6f",x"4c",x"87",x"c1"),
  1055 => (x"6e",x"69",x"64",x"61"),
  1056 => (x"2e",x"2e",x"2e",x"67"),
  1057 => (x"1e",x"73",x"1e",x"00"),
  1058 => (x"c2",x"49",x"4a",x"71"),
  1059 => (x"81",x"bf",x"d8",x"ea"),
  1060 => (x"87",x"ef",x"fb",x"71"),
  1061 => (x"02",x"9b",x"4b",x"70"),
  1062 => (x"e7",x"49",x"87",x"c4"),
  1063 => (x"ea",x"c2",x"87",x"e9"),
  1064 => (x"78",x"c0",x"48",x"d8"),
  1065 => (x"d7",x"dd",x"49",x"c1"),
  1066 => (x"87",x"d3",x"fb",x"87"),
  1067 => (x"c1",x"49",x"c0",x"1e"),
  1068 => (x"26",x"87",x"e3",x"c0"),
  1069 => (x"4a",x"71",x"1e",x"4f"),
  1070 => (x"c1",x"91",x"cb",x"49"),
  1071 => (x"c8",x"81",x"d4",x"e3"),
  1072 => (x"c2",x"48",x"11",x"81"),
  1073 => (x"c2",x"58",x"c4",x"ea"),
  1074 => (x"c0",x"48",x"d8",x"ea"),
  1075 => (x"dc",x"49",x"c1",x"78"),
  1076 => (x"4f",x"26",x"87",x"ee"),
  1077 => (x"02",x"99",x"71",x"1e"),
  1078 => (x"e4",x"c1",x"87",x"d2"),
  1079 => (x"50",x"c0",x"48",x"e9"),
  1080 => (x"c2",x"c1",x"80",x"f7"),
  1081 => (x"e3",x"c1",x"40",x"f5"),
  1082 => (x"87",x"ce",x"78",x"cd"),
  1083 => (x"48",x"e5",x"e4",x"c1"),
  1084 => (x"78",x"c6",x"e3",x"c1"),
  1085 => (x"c2",x"c1",x"80",x"fc"),
  1086 => (x"4f",x"26",x"78",x"ec"),
  1087 => (x"5c",x"5b",x"5e",x"0e"),
  1088 => (x"86",x"f4",x"0e",x"5d"),
  1089 => (x"4d",x"ce",x"dd",x"c2"),
  1090 => (x"a6",x"c4",x"4c",x"c0"),
  1091 => (x"c2",x"78",x"c0",x"48"),
  1092 => (x"48",x"bf",x"d8",x"ea"),
  1093 => (x"c1",x"06",x"a8",x"c0"),
  1094 => (x"dd",x"c2",x"87",x"c0"),
  1095 => (x"02",x"98",x"48",x"ce"),
  1096 => (x"c0",x"87",x"f7",x"c0"),
  1097 => (x"c8",x"1e",x"cf",x"f6"),
  1098 => (x"87",x"c7",x"02",x"66"),
  1099 => (x"c0",x"48",x"a6",x"c4"),
  1100 => (x"c4",x"87",x"c5",x"78"),
  1101 => (x"78",x"c1",x"48",x"a6"),
  1102 => (x"e6",x"49",x"66",x"c4"),
  1103 => (x"86",x"c4",x"87",x"c0"),
  1104 => (x"84",x"c1",x"4d",x"70"),
  1105 => (x"c1",x"48",x"66",x"c4"),
  1106 => (x"58",x"a6",x"c8",x"80"),
  1107 => (x"bf",x"d8",x"ea",x"c2"),
  1108 => (x"87",x"c6",x"03",x"ac"),
  1109 => (x"ff",x"05",x"9d",x"75"),
  1110 => (x"4c",x"c0",x"87",x"c9"),
  1111 => (x"c3",x"02",x"9d",x"75"),
  1112 => (x"f6",x"c0",x"87",x"dc"),
  1113 => (x"66",x"c8",x"1e",x"cf"),
  1114 => (x"cc",x"87",x"c7",x"02"),
  1115 => (x"78",x"c0",x"48",x"a6"),
  1116 => (x"a6",x"cc",x"87",x"c5"),
  1117 => (x"cc",x"78",x"c1",x"48"),
  1118 => (x"c1",x"e5",x"49",x"66"),
  1119 => (x"70",x"86",x"c4",x"87"),
  1120 => (x"02",x"98",x"48",x"7e"),
  1121 => (x"49",x"87",x"e4",x"c2"),
  1122 => (x"69",x"97",x"81",x"cb"),
  1123 => (x"02",x"99",x"d0",x"49"),
  1124 => (x"74",x"87",x"d4",x"c1"),
  1125 => (x"c1",x"91",x"cb",x"49"),
  1126 => (x"c1",x"81",x"d4",x"e3"),
  1127 => (x"c8",x"79",x"c5",x"c2"),
  1128 => (x"51",x"ff",x"c3",x"81"),
  1129 => (x"91",x"de",x"49",x"74"),
  1130 => (x"4d",x"ec",x"ea",x"c2"),
  1131 => (x"c1",x"c2",x"85",x"71"),
  1132 => (x"a5",x"c1",x"7d",x"97"),
  1133 => (x"51",x"e0",x"c0",x"49"),
  1134 => (x"97",x"de",x"e5",x"c2"),
  1135 => (x"87",x"d2",x"02",x"bf"),
  1136 => (x"a5",x"c2",x"84",x"c1"),
  1137 => (x"de",x"e5",x"c2",x"4b"),
  1138 => (x"fe",x"49",x"db",x"4a"),
  1139 => (x"c1",x"87",x"d8",x"fb"),
  1140 => (x"a5",x"cd",x"87",x"d9"),
  1141 => (x"c1",x"51",x"c0",x"49"),
  1142 => (x"4b",x"a5",x"c2",x"84"),
  1143 => (x"49",x"cb",x"4a",x"6e"),
  1144 => (x"87",x"c3",x"fb",x"fe"),
  1145 => (x"74",x"87",x"c4",x"c1"),
  1146 => (x"c1",x"91",x"cb",x"49"),
  1147 => (x"c1",x"81",x"d4",x"e3"),
  1148 => (x"c2",x"79",x"c2",x"c0"),
  1149 => (x"bf",x"97",x"de",x"e5"),
  1150 => (x"74",x"87",x"d8",x"02"),
  1151 => (x"c1",x"91",x"de",x"49"),
  1152 => (x"ec",x"ea",x"c2",x"84"),
  1153 => (x"c2",x"83",x"71",x"4b"),
  1154 => (x"dd",x"4a",x"de",x"e5"),
  1155 => (x"d6",x"fa",x"fe",x"49"),
  1156 => (x"74",x"87",x"d8",x"87"),
  1157 => (x"c2",x"93",x"de",x"4b"),
  1158 => (x"cb",x"83",x"ec",x"ea"),
  1159 => (x"51",x"c0",x"49",x"a3"),
  1160 => (x"6e",x"73",x"84",x"c1"),
  1161 => (x"fe",x"49",x"cb",x"4a"),
  1162 => (x"c4",x"87",x"fc",x"f9"),
  1163 => (x"80",x"c1",x"48",x"66"),
  1164 => (x"c7",x"58",x"a6",x"c8"),
  1165 => (x"c5",x"c0",x"03",x"ac"),
  1166 => (x"fc",x"05",x"6e",x"87"),
  1167 => (x"48",x"74",x"87",x"e4"),
  1168 => (x"f6",x"f4",x"8e",x"f4"),
  1169 => (x"1e",x"73",x"1e",x"87"),
  1170 => (x"cb",x"49",x"4b",x"71"),
  1171 => (x"d4",x"e3",x"c1",x"91"),
  1172 => (x"4a",x"a1",x"c8",x"81"),
  1173 => (x"48",x"c0",x"e3",x"c1"),
  1174 => (x"a1",x"c9",x"50",x"12"),
  1175 => (x"ee",x"f8",x"c0",x"4a"),
  1176 => (x"ca",x"50",x"12",x"48"),
  1177 => (x"c1",x"e3",x"c1",x"81"),
  1178 => (x"c1",x"50",x"11",x"48"),
  1179 => (x"bf",x"97",x"c1",x"e3"),
  1180 => (x"49",x"c0",x"1e",x"49"),
  1181 => (x"c2",x"87",x"cb",x"f5"),
  1182 => (x"de",x"48",x"c0",x"ea"),
  1183 => (x"d5",x"49",x"c1",x"78"),
  1184 => (x"f3",x"26",x"87",x"fe"),
  1185 => (x"5e",x"0e",x"87",x"f9"),
  1186 => (x"0e",x"5d",x"5c",x"5b"),
  1187 => (x"4d",x"71",x"86",x"f4"),
  1188 => (x"c1",x"91",x"cb",x"49"),
  1189 => (x"c8",x"81",x"d4",x"e3"),
  1190 => (x"a1",x"ca",x"4a",x"a1"),
  1191 => (x"48",x"a6",x"c4",x"7e"),
  1192 => (x"bf",x"c8",x"ee",x"c2"),
  1193 => (x"bf",x"97",x"6e",x"78"),
  1194 => (x"4c",x"66",x"c4",x"4b"),
  1195 => (x"48",x"12",x"2c",x"73"),
  1196 => (x"70",x"58",x"a6",x"cc"),
  1197 => (x"c9",x"84",x"c1",x"9c"),
  1198 => (x"49",x"69",x"97",x"81"),
  1199 => (x"c2",x"04",x"ac",x"b7"),
  1200 => (x"6e",x"4c",x"c0",x"87"),
  1201 => (x"c8",x"4a",x"bf",x"97"),
  1202 => (x"31",x"72",x"49",x"66"),
  1203 => (x"66",x"c4",x"b9",x"ff"),
  1204 => (x"72",x"48",x"74",x"99"),
  1205 => (x"48",x"4a",x"70",x"30"),
  1206 => (x"ee",x"c2",x"b0",x"71"),
  1207 => (x"e4",x"c0",x"58",x"cc"),
  1208 => (x"49",x"c0",x"87",x"cf"),
  1209 => (x"75",x"87",x"d9",x"d4"),
  1210 => (x"c4",x"f6",x"c0",x"49"),
  1211 => (x"f2",x"8e",x"f4",x"87"),
  1212 => (x"73",x"1e",x"87",x"c9"),
  1213 => (x"49",x"4b",x"71",x"1e"),
  1214 => (x"73",x"87",x"cb",x"fe"),
  1215 => (x"87",x"c6",x"fe",x"49"),
  1216 => (x"1e",x"87",x"fc",x"f1"),
  1217 => (x"4b",x"71",x"1e",x"73"),
  1218 => (x"02",x"4a",x"a3",x"c6"),
  1219 => (x"c1",x"87",x"e3",x"c0"),
  1220 => (x"87",x"d6",x"02",x"8a"),
  1221 => (x"e8",x"c1",x"02",x"8a"),
  1222 => (x"c1",x"02",x"8a",x"87"),
  1223 => (x"02",x"8a",x"87",x"ca"),
  1224 => (x"8a",x"87",x"ef",x"c0"),
  1225 => (x"c1",x"87",x"d9",x"02"),
  1226 => (x"49",x"c7",x"87",x"e9"),
  1227 => (x"c1",x"87",x"c6",x"f6"),
  1228 => (x"ea",x"c2",x"87",x"ec"),
  1229 => (x"78",x"df",x"48",x"c0"),
  1230 => (x"c3",x"d3",x"49",x"c1"),
  1231 => (x"87",x"de",x"c1",x"87"),
  1232 => (x"bf",x"d8",x"ea",x"c2"),
  1233 => (x"87",x"cb",x"c1",x"02"),
  1234 => (x"c2",x"88",x"c1",x"48"),
  1235 => (x"c1",x"58",x"dc",x"ea"),
  1236 => (x"ea",x"c2",x"87",x"c1"),
  1237 => (x"c0",x"02",x"bf",x"dc"),
  1238 => (x"ea",x"c2",x"87",x"f9"),
  1239 => (x"c1",x"48",x"bf",x"d8"),
  1240 => (x"dc",x"ea",x"c2",x"80"),
  1241 => (x"87",x"eb",x"c0",x"58"),
  1242 => (x"bf",x"d8",x"ea",x"c2"),
  1243 => (x"c2",x"89",x"c6",x"49"),
  1244 => (x"c0",x"59",x"dc",x"ea"),
  1245 => (x"da",x"03",x"a9",x"b7"),
  1246 => (x"d8",x"ea",x"c2",x"87"),
  1247 => (x"d2",x"78",x"c0",x"48"),
  1248 => (x"dc",x"ea",x"c2",x"87"),
  1249 => (x"87",x"cb",x"02",x"bf"),
  1250 => (x"bf",x"d8",x"ea",x"c2"),
  1251 => (x"c2",x"80",x"c6",x"48"),
  1252 => (x"c0",x"58",x"dc",x"ea"),
  1253 => (x"87",x"e8",x"d1",x"49"),
  1254 => (x"f3",x"c0",x"49",x"73"),
  1255 => (x"de",x"ef",x"87",x"d3"),
  1256 => (x"5b",x"5e",x"0e",x"87"),
  1257 => (x"ff",x"0e",x"5d",x"5c"),
  1258 => (x"a6",x"dc",x"86",x"d4"),
  1259 => (x"48",x"a6",x"c8",x"59"),
  1260 => (x"80",x"c4",x"78",x"c0"),
  1261 => (x"78",x"66",x"c0",x"c1"),
  1262 => (x"78",x"c1",x"80",x"c4"),
  1263 => (x"78",x"c1",x"80",x"c4"),
  1264 => (x"48",x"dc",x"ea",x"c2"),
  1265 => (x"ea",x"c2",x"78",x"c1"),
  1266 => (x"de",x"48",x"bf",x"c0"),
  1267 => (x"87",x"c9",x"05",x"a8"),
  1268 => (x"cc",x"87",x"e9",x"f4"),
  1269 => (x"e6",x"cf",x"58",x"a6"),
  1270 => (x"87",x"e2",x"e3",x"87"),
  1271 => (x"e3",x"87",x"c4",x"e4"),
  1272 => (x"4c",x"70",x"87",x"d1"),
  1273 => (x"02",x"ac",x"fb",x"c0"),
  1274 => (x"d8",x"87",x"fb",x"c1"),
  1275 => (x"ed",x"c1",x"05",x"66"),
  1276 => (x"66",x"fc",x"c0",x"87"),
  1277 => (x"6a",x"82",x"c4",x"4a"),
  1278 => (x"c1",x"1e",x"72",x"7e"),
  1279 => (x"c4",x"48",x"f4",x"df"),
  1280 => (x"a1",x"c8",x"49",x"66"),
  1281 => (x"71",x"41",x"20",x"4a"),
  1282 => (x"87",x"f9",x"05",x"aa"),
  1283 => (x"4a",x"26",x"51",x"10"),
  1284 => (x"48",x"66",x"fc",x"c0"),
  1285 => (x"78",x"c5",x"c9",x"c1"),
  1286 => (x"81",x"c7",x"49",x"6a"),
  1287 => (x"fc",x"c0",x"51",x"74"),
  1288 => (x"81",x"c8",x"49",x"66"),
  1289 => (x"fc",x"c0",x"51",x"c1"),
  1290 => (x"81",x"c9",x"49",x"66"),
  1291 => (x"fc",x"c0",x"51",x"c0"),
  1292 => (x"81",x"ca",x"49",x"66"),
  1293 => (x"1e",x"c1",x"51",x"c0"),
  1294 => (x"49",x"6a",x"1e",x"d8"),
  1295 => (x"f6",x"e2",x"81",x"c8"),
  1296 => (x"c1",x"86",x"c8",x"87"),
  1297 => (x"c0",x"48",x"66",x"c0"),
  1298 => (x"87",x"c7",x"01",x"a8"),
  1299 => (x"c1",x"48",x"a6",x"c8"),
  1300 => (x"c1",x"87",x"ce",x"78"),
  1301 => (x"c1",x"48",x"66",x"c0"),
  1302 => (x"58",x"a6",x"d0",x"88"),
  1303 => (x"c2",x"e2",x"87",x"c3"),
  1304 => (x"48",x"a6",x"d0",x"87"),
  1305 => (x"9c",x"74",x"78",x"c2"),
  1306 => (x"87",x"cf",x"cd",x"02"),
  1307 => (x"c1",x"48",x"66",x"c8"),
  1308 => (x"03",x"a8",x"66",x"c4"),
  1309 => (x"dc",x"87",x"c4",x"cd"),
  1310 => (x"78",x"c0",x"48",x"a6"),
  1311 => (x"78",x"c0",x"80",x"e8"),
  1312 => (x"70",x"87",x"f0",x"e0"),
  1313 => (x"ac",x"d0",x"c1",x"4c"),
  1314 => (x"87",x"d7",x"c2",x"05"),
  1315 => (x"e3",x"7e",x"66",x"c4"),
  1316 => (x"a6",x"c8",x"87",x"d4"),
  1317 => (x"87",x"db",x"e0",x"58"),
  1318 => (x"ec",x"c0",x"4c",x"70"),
  1319 => (x"ed",x"c1",x"05",x"ac"),
  1320 => (x"49",x"66",x"c8",x"87"),
  1321 => (x"fc",x"c0",x"91",x"cb"),
  1322 => (x"a1",x"c4",x"81",x"66"),
  1323 => (x"c8",x"4d",x"6a",x"4a"),
  1324 => (x"66",x"c4",x"4a",x"a1"),
  1325 => (x"f5",x"c2",x"c1",x"52"),
  1326 => (x"f6",x"df",x"ff",x"79"),
  1327 => (x"9c",x"4c",x"70",x"87"),
  1328 => (x"c0",x"87",x"d9",x"02"),
  1329 => (x"d3",x"02",x"ac",x"fb"),
  1330 => (x"ff",x"55",x"74",x"87"),
  1331 => (x"70",x"87",x"e4",x"df"),
  1332 => (x"c7",x"02",x"9c",x"4c"),
  1333 => (x"ac",x"fb",x"c0",x"87"),
  1334 => (x"87",x"ed",x"ff",x"05"),
  1335 => (x"c2",x"55",x"e0",x"c0"),
  1336 => (x"97",x"c0",x"55",x"c1"),
  1337 => (x"48",x"66",x"d8",x"7d"),
  1338 => (x"db",x"05",x"a8",x"6e"),
  1339 => (x"48",x"66",x"c8",x"87"),
  1340 => (x"04",x"a8",x"66",x"cc"),
  1341 => (x"66",x"c8",x"87",x"ca"),
  1342 => (x"cc",x"80",x"c1",x"48"),
  1343 => (x"87",x"c8",x"58",x"a6"),
  1344 => (x"c1",x"48",x"66",x"cc"),
  1345 => (x"58",x"a6",x"d0",x"88"),
  1346 => (x"87",x"e7",x"de",x"ff"),
  1347 => (x"d0",x"c1",x"4c",x"70"),
  1348 => (x"87",x"c8",x"05",x"ac"),
  1349 => (x"c1",x"48",x"66",x"d4"),
  1350 => (x"58",x"a6",x"d8",x"80"),
  1351 => (x"02",x"ac",x"d0",x"c1"),
  1352 => (x"c4",x"87",x"e9",x"fd"),
  1353 => (x"66",x"d8",x"48",x"66"),
  1354 => (x"e0",x"c9",x"05",x"a8"),
  1355 => (x"a6",x"e0",x"c0",x"87"),
  1356 => (x"74",x"78",x"c0",x"48"),
  1357 => (x"88",x"fb",x"c0",x"48"),
  1358 => (x"98",x"48",x"7e",x"70"),
  1359 => (x"87",x"e2",x"c9",x"02"),
  1360 => (x"70",x"88",x"cb",x"48"),
  1361 => (x"02",x"98",x"48",x"7e"),
  1362 => (x"48",x"87",x"cd",x"c1"),
  1363 => (x"7e",x"70",x"88",x"c9"),
  1364 => (x"c3",x"02",x"98",x"48"),
  1365 => (x"c4",x"48",x"87",x"fe"),
  1366 => (x"48",x"7e",x"70",x"88"),
  1367 => (x"87",x"ce",x"02",x"98"),
  1368 => (x"70",x"88",x"c1",x"48"),
  1369 => (x"02",x"98",x"48",x"7e"),
  1370 => (x"c8",x"87",x"e9",x"c3"),
  1371 => (x"a6",x"dc",x"87",x"d6"),
  1372 => (x"78",x"f0",x"c0",x"48"),
  1373 => (x"87",x"fb",x"dc",x"ff"),
  1374 => (x"ec",x"c0",x"4c",x"70"),
  1375 => (x"c4",x"c0",x"02",x"ac"),
  1376 => (x"a6",x"e0",x"c0",x"87"),
  1377 => (x"ac",x"ec",x"c0",x"5c"),
  1378 => (x"ff",x"87",x"cd",x"02"),
  1379 => (x"70",x"87",x"e4",x"dc"),
  1380 => (x"ac",x"ec",x"c0",x"4c"),
  1381 => (x"87",x"f3",x"ff",x"05"),
  1382 => (x"02",x"ac",x"ec",x"c0"),
  1383 => (x"ff",x"87",x"c4",x"c0"),
  1384 => (x"c0",x"87",x"d0",x"dc"),
  1385 => (x"d0",x"1e",x"ca",x"1e"),
  1386 => (x"91",x"cb",x"49",x"66"),
  1387 => (x"48",x"66",x"c4",x"c1"),
  1388 => (x"a6",x"cc",x"80",x"71"),
  1389 => (x"48",x"66",x"c8",x"58"),
  1390 => (x"a6",x"d0",x"80",x"c4"),
  1391 => (x"bf",x"66",x"cc",x"58"),
  1392 => (x"f2",x"dc",x"ff",x"49"),
  1393 => (x"de",x"1e",x"c1",x"87"),
  1394 => (x"bf",x"66",x"d4",x"1e"),
  1395 => (x"e6",x"dc",x"ff",x"49"),
  1396 => (x"70",x"86",x"d0",x"87"),
  1397 => (x"08",x"c0",x"48",x"49"),
  1398 => (x"a6",x"e8",x"c0",x"88"),
  1399 => (x"06",x"a8",x"c0",x"58"),
  1400 => (x"c0",x"87",x"ee",x"c0"),
  1401 => (x"dd",x"48",x"66",x"e4"),
  1402 => (x"e4",x"c0",x"03",x"a8"),
  1403 => (x"bf",x"66",x"c4",x"87"),
  1404 => (x"66",x"e4",x"c0",x"49"),
  1405 => (x"51",x"e0",x"c0",x"81"),
  1406 => (x"49",x"66",x"e4",x"c0"),
  1407 => (x"66",x"c4",x"81",x"c1"),
  1408 => (x"c1",x"c2",x"81",x"bf"),
  1409 => (x"66",x"e4",x"c0",x"51"),
  1410 => (x"c4",x"81",x"c2",x"49"),
  1411 => (x"c0",x"81",x"bf",x"66"),
  1412 => (x"c1",x"48",x"6e",x"51"),
  1413 => (x"6e",x"78",x"c5",x"c9"),
  1414 => (x"d0",x"81",x"c8",x"49"),
  1415 => (x"49",x"6e",x"51",x"66"),
  1416 => (x"66",x"d4",x"81",x"c9"),
  1417 => (x"ca",x"49",x"6e",x"51"),
  1418 => (x"51",x"66",x"dc",x"81"),
  1419 => (x"c1",x"48",x"66",x"d0"),
  1420 => (x"58",x"a6",x"d4",x"80"),
  1421 => (x"cc",x"48",x"66",x"c8"),
  1422 => (x"c0",x"04",x"a8",x"66"),
  1423 => (x"66",x"c8",x"87",x"cb"),
  1424 => (x"cc",x"80",x"c1",x"48"),
  1425 => (x"d9",x"c5",x"58",x"a6"),
  1426 => (x"48",x"66",x"cc",x"87"),
  1427 => (x"a6",x"d0",x"88",x"c1"),
  1428 => (x"87",x"ce",x"c5",x"58"),
  1429 => (x"87",x"ce",x"dc",x"ff"),
  1430 => (x"58",x"a6",x"e8",x"c0"),
  1431 => (x"87",x"c6",x"dc",x"ff"),
  1432 => (x"58",x"a6",x"e0",x"c0"),
  1433 => (x"05",x"a8",x"ec",x"c0"),
  1434 => (x"dc",x"87",x"ca",x"c0"),
  1435 => (x"e4",x"c0",x"48",x"a6"),
  1436 => (x"c4",x"c0",x"78",x"66"),
  1437 => (x"fa",x"d8",x"ff",x"87"),
  1438 => (x"49",x"66",x"c8",x"87"),
  1439 => (x"fc",x"c0",x"91",x"cb"),
  1440 => (x"80",x"71",x"48",x"66"),
  1441 => (x"c8",x"4a",x"7e",x"70"),
  1442 => (x"ca",x"49",x"6e",x"82"),
  1443 => (x"66",x"e4",x"c0",x"81"),
  1444 => (x"49",x"66",x"dc",x"51"),
  1445 => (x"e4",x"c0",x"81",x"c1"),
  1446 => (x"48",x"c1",x"89",x"66"),
  1447 => (x"49",x"70",x"30",x"71"),
  1448 => (x"97",x"71",x"89",x"c1"),
  1449 => (x"c8",x"ee",x"c2",x"7a"),
  1450 => (x"e4",x"c0",x"49",x"bf"),
  1451 => (x"6a",x"97",x"29",x"66"),
  1452 => (x"98",x"71",x"48",x"4a"),
  1453 => (x"58",x"a6",x"ec",x"c0"),
  1454 => (x"81",x"c4",x"49",x"6e"),
  1455 => (x"66",x"d8",x"4d",x"69"),
  1456 => (x"a8",x"66",x"c4",x"48"),
  1457 => (x"87",x"c8",x"c0",x"02"),
  1458 => (x"c0",x"48",x"a6",x"c4"),
  1459 => (x"87",x"c5",x"c0",x"78"),
  1460 => (x"c1",x"48",x"a6",x"c4"),
  1461 => (x"1e",x"66",x"c4",x"78"),
  1462 => (x"75",x"1e",x"e0",x"c0"),
  1463 => (x"d6",x"d8",x"ff",x"49"),
  1464 => (x"70",x"86",x"c8",x"87"),
  1465 => (x"ac",x"b7",x"c0",x"4c"),
  1466 => (x"87",x"d4",x"c1",x"06"),
  1467 => (x"e0",x"c0",x"85",x"74"),
  1468 => (x"75",x"89",x"74",x"49"),
  1469 => (x"fd",x"df",x"c1",x"4b"),
  1470 => (x"e6",x"fe",x"71",x"4a"),
  1471 => (x"85",x"c2",x"87",x"e9"),
  1472 => (x"48",x"66",x"e0",x"c0"),
  1473 => (x"e4",x"c0",x"80",x"c1"),
  1474 => (x"e8",x"c0",x"58",x"a6"),
  1475 => (x"81",x"c1",x"49",x"66"),
  1476 => (x"c0",x"02",x"a9",x"70"),
  1477 => (x"a6",x"c4",x"87",x"c8"),
  1478 => (x"c0",x"78",x"c0",x"48"),
  1479 => (x"a6",x"c4",x"87",x"c5"),
  1480 => (x"c4",x"78",x"c1",x"48"),
  1481 => (x"a4",x"c2",x"1e",x"66"),
  1482 => (x"48",x"e0",x"c0",x"49"),
  1483 => (x"49",x"70",x"88",x"71"),
  1484 => (x"ff",x"49",x"75",x"1e"),
  1485 => (x"c8",x"87",x"c0",x"d7"),
  1486 => (x"a8",x"b7",x"c0",x"86"),
  1487 => (x"87",x"c0",x"ff",x"01"),
  1488 => (x"02",x"66",x"e0",x"c0"),
  1489 => (x"6e",x"87",x"d1",x"c0"),
  1490 => (x"c0",x"81",x"c9",x"49"),
  1491 => (x"6e",x"51",x"66",x"e0"),
  1492 => (x"c6",x"ca",x"c1",x"48"),
  1493 => (x"87",x"cc",x"c0",x"78"),
  1494 => (x"81",x"c9",x"49",x"6e"),
  1495 => (x"48",x"6e",x"51",x"c2"),
  1496 => (x"78",x"f2",x"cb",x"c1"),
  1497 => (x"cc",x"48",x"66",x"c8"),
  1498 => (x"c0",x"04",x"a8",x"66"),
  1499 => (x"66",x"c8",x"87",x"cb"),
  1500 => (x"cc",x"80",x"c1",x"48"),
  1501 => (x"e9",x"c0",x"58",x"a6"),
  1502 => (x"48",x"66",x"cc",x"87"),
  1503 => (x"a6",x"d0",x"88",x"c1"),
  1504 => (x"87",x"de",x"c0",x"58"),
  1505 => (x"87",x"db",x"d5",x"ff"),
  1506 => (x"d5",x"c0",x"4c",x"70"),
  1507 => (x"ac",x"c6",x"c1",x"87"),
  1508 => (x"87",x"c8",x"c0",x"05"),
  1509 => (x"c1",x"48",x"66",x"d0"),
  1510 => (x"58",x"a6",x"d4",x"80"),
  1511 => (x"87",x"c3",x"d5",x"ff"),
  1512 => (x"66",x"d4",x"4c",x"70"),
  1513 => (x"d8",x"80",x"c1",x"48"),
  1514 => (x"9c",x"74",x"58",x"a6"),
  1515 => (x"87",x"cb",x"c0",x"02"),
  1516 => (x"c1",x"48",x"66",x"c8"),
  1517 => (x"04",x"a8",x"66",x"c4"),
  1518 => (x"ff",x"87",x"fc",x"f2"),
  1519 => (x"c8",x"87",x"db",x"d4"),
  1520 => (x"a8",x"c7",x"48",x"66"),
  1521 => (x"87",x"e5",x"c0",x"03"),
  1522 => (x"48",x"dc",x"ea",x"c2"),
  1523 => (x"66",x"c8",x"78",x"c0"),
  1524 => (x"c0",x"91",x"cb",x"49"),
  1525 => (x"c4",x"81",x"66",x"fc"),
  1526 => (x"4a",x"6a",x"4a",x"a1"),
  1527 => (x"c8",x"79",x"52",x"c0"),
  1528 => (x"80",x"c1",x"48",x"66"),
  1529 => (x"c7",x"58",x"a6",x"cc"),
  1530 => (x"db",x"ff",x"04",x"a8"),
  1531 => (x"8e",x"d4",x"ff",x"87"),
  1532 => (x"87",x"c7",x"de",x"ff"),
  1533 => (x"64",x"61",x"6f",x"4c"),
  1534 => (x"20",x"2e",x"2a",x"20"),
  1535 => (x"00",x"20",x"3a",x"00"),
  1536 => (x"71",x"1e",x"73",x"1e"),
  1537 => (x"c6",x"02",x"9b",x"4b"),
  1538 => (x"d8",x"ea",x"c2",x"87"),
  1539 => (x"c7",x"78",x"c0",x"48"),
  1540 => (x"d8",x"ea",x"c2",x"1e"),
  1541 => (x"e3",x"c1",x"1e",x"bf"),
  1542 => (x"ea",x"c2",x"1e",x"d4"),
  1543 => (x"ed",x"49",x"bf",x"c0"),
  1544 => (x"86",x"cc",x"87",x"ff"),
  1545 => (x"bf",x"c0",x"ea",x"c2"),
  1546 => (x"87",x"e8",x"e2",x"49"),
  1547 => (x"c8",x"02",x"9b",x"73"),
  1548 => (x"d4",x"e3",x"c1",x"87"),
  1549 => (x"ca",x"e2",x"c0",x"49"),
  1550 => (x"c2",x"dd",x"ff",x"87"),
  1551 => (x"ca",x"c7",x"1e",x"87"),
  1552 => (x"fe",x"49",x"c1",x"87"),
  1553 => (x"ea",x"c2",x"87",x"fa"),
  1554 => (x"50",x"c0",x"48",x"e0"),
  1555 => (x"87",x"c7",x"ea",x"fe"),
  1556 => (x"cd",x"02",x"98",x"70"),
  1557 => (x"c1",x"f3",x"fe",x"87"),
  1558 => (x"02",x"98",x"70",x"87"),
  1559 => (x"4a",x"c1",x"87",x"c4"),
  1560 => (x"4a",x"c0",x"87",x"c2"),
  1561 => (x"ce",x"05",x"9a",x"72"),
  1562 => (x"c1",x"1e",x"c0",x"87"),
  1563 => (x"c0",x"49",x"ea",x"e2"),
  1564 => (x"c4",x"87",x"fb",x"ef"),
  1565 => (x"c2",x"87",x"fe",x"86"),
  1566 => (x"c0",x"48",x"d8",x"ea"),
  1567 => (x"c0",x"ea",x"c2",x"78"),
  1568 => (x"1e",x"78",x"c0",x"48"),
  1569 => (x"49",x"f5",x"e2",x"c1"),
  1570 => (x"87",x"e2",x"ef",x"c0"),
  1571 => (x"f8",x"c0",x"1e",x"c0"),
  1572 => (x"49",x"70",x"87",x"f4"),
  1573 => (x"87",x"d6",x"ef",x"c0"),
  1574 => (x"ed",x"c2",x"86",x"c8"),
  1575 => (x"df",x"e2",x"c0",x"87"),
  1576 => (x"d4",x"f3",x"c0",x"87"),
  1577 => (x"87",x"f5",x"ff",x"87"),
  1578 => (x"44",x"53",x"4f",x"26"),
  1579 => (x"69",x"61",x"66",x"20"),
  1580 => (x"2e",x"64",x"65",x"6c"),
  1581 => (x"6f",x"6f",x"42",x"00"),
  1582 => (x"67",x"6e",x"69",x"74"),
  1583 => (x"00",x"2e",x"2e",x"2e"),
  1584 => (x"00",x"01",x"00",x"00"),
  1585 => (x"20",x"80",x"00",x"00"),
  1586 => (x"74",x"69",x"78",x"45"),
  1587 => (x"42",x"20",x"80",x"00"),
  1588 => (x"00",x"6b",x"63",x"61"),
  1589 => (x"00",x"00",x"10",x"02"),
  1590 => (x"00",x"00",x"2a",x"ac"),
  1591 => (x"02",x"00",x"00",x"00"),
  1592 => (x"ca",x"00",x"00",x"10"),
  1593 => (x"00",x"00",x"00",x"2a"),
  1594 => (x"10",x"02",x"00",x"00"),
  1595 => (x"2a",x"e8",x"00",x"00"),
  1596 => (x"00",x"00",x"00",x"00"),
  1597 => (x"00",x"10",x"02",x"00"),
  1598 => (x"00",x"2b",x"06",x"00"),
  1599 => (x"00",x"00",x"00",x"00"),
  1600 => (x"00",x"00",x"10",x"02"),
  1601 => (x"00",x"00",x"2b",x"24"),
  1602 => (x"02",x"00",x"00",x"00"),
  1603 => (x"42",x"00",x"00",x"10"),
  1604 => (x"00",x"00",x"00",x"2b"),
  1605 => (x"10",x"02",x"00",x"00"),
  1606 => (x"2b",x"60",x"00",x"00"),
  1607 => (x"00",x"00",x"00",x"00"),
  1608 => (x"00",x"10",x"b5",x"00"),
  1609 => (x"00",x"00",x"00",x"00"),
  1610 => (x"00",x"00",x"00",x"00"),
  1611 => (x"00",x"00",x"13",x"03"),
  1612 => (x"00",x"00",x"00",x"00"),
  1613 => (x"1e",x"00",x"00",x"00"),
  1614 => (x"c0",x"48",x"f0",x"fe"),
  1615 => (x"79",x"09",x"cd",x"78"),
  1616 => (x"1e",x"4f",x"26",x"09"),
  1617 => (x"48",x"bf",x"f0",x"fe"),
  1618 => (x"fe",x"1e",x"4f",x"26"),
  1619 => (x"78",x"c1",x"48",x"f0"),
  1620 => (x"fe",x"1e",x"4f",x"26"),
  1621 => (x"78",x"c0",x"48",x"f0"),
  1622 => (x"71",x"1e",x"4f",x"26"),
  1623 => (x"51",x"52",x"c0",x"4a"),
  1624 => (x"5e",x"0e",x"4f",x"26"),
  1625 => (x"0e",x"5d",x"5c",x"5b"),
  1626 => (x"4d",x"71",x"86",x"f4"),
  1627 => (x"c1",x"7e",x"6d",x"97"),
  1628 => (x"6c",x"97",x"4c",x"a5"),
  1629 => (x"58",x"a6",x"c8",x"48"),
  1630 => (x"66",x"c4",x"48",x"6e"),
  1631 => (x"87",x"c5",x"05",x"a8"),
  1632 => (x"e6",x"c0",x"48",x"ff"),
  1633 => (x"87",x"ca",x"ff",x"87"),
  1634 => (x"97",x"49",x"a5",x"c2"),
  1635 => (x"a3",x"71",x"4b",x"6c"),
  1636 => (x"4b",x"6b",x"97",x"4b"),
  1637 => (x"6e",x"7e",x"6c",x"97"),
  1638 => (x"c8",x"80",x"c1",x"48"),
  1639 => (x"98",x"c7",x"58",x"a6"),
  1640 => (x"70",x"58",x"a6",x"cc"),
  1641 => (x"e1",x"fe",x"7c",x"97"),
  1642 => (x"f4",x"48",x"73",x"87"),
  1643 => (x"26",x"4d",x"26",x"8e"),
  1644 => (x"26",x"4b",x"26",x"4c"),
  1645 => (x"5b",x"5e",x"0e",x"4f"),
  1646 => (x"86",x"f4",x"0e",x"5c"),
  1647 => (x"66",x"d8",x"4c",x"71"),
  1648 => (x"9a",x"ff",x"c3",x"4a"),
  1649 => (x"97",x"4b",x"a4",x"c2"),
  1650 => (x"a1",x"73",x"49",x"6c"),
  1651 => (x"97",x"51",x"72",x"49"),
  1652 => (x"48",x"6e",x"7e",x"6c"),
  1653 => (x"a6",x"c8",x"80",x"c1"),
  1654 => (x"cc",x"98",x"c7",x"58"),
  1655 => (x"54",x"70",x"58",x"a6"),
  1656 => (x"ca",x"ff",x"8e",x"f4"),
  1657 => (x"fd",x"1e",x"1e",x"87"),
  1658 => (x"bf",x"e0",x"87",x"e8"),
  1659 => (x"e0",x"c0",x"49",x"4a"),
  1660 => (x"cb",x"02",x"99",x"c0"),
  1661 => (x"c2",x"1e",x"72",x"87"),
  1662 => (x"fe",x"49",x"fe",x"ed"),
  1663 => (x"86",x"c4",x"87",x"f7"),
  1664 => (x"70",x"87",x"c0",x"fd"),
  1665 => (x"87",x"c2",x"fd",x"7e"),
  1666 => (x"1e",x"4f",x"26",x"26"),
  1667 => (x"49",x"fe",x"ed",x"c2"),
  1668 => (x"c1",x"87",x"c7",x"fd"),
  1669 => (x"fc",x"49",x"e5",x"e7"),
  1670 => (x"ee",x"c3",x"87",x"dd"),
  1671 => (x"0e",x"4f",x"26",x"87"),
  1672 => (x"5d",x"5c",x"5b",x"5e"),
  1673 => (x"c2",x"4d",x"71",x"0e"),
  1674 => (x"fc",x"49",x"fe",x"ed"),
  1675 => (x"4b",x"70",x"87",x"f4"),
  1676 => (x"04",x"ab",x"b7",x"c0"),
  1677 => (x"c3",x"87",x"c2",x"c3"),
  1678 => (x"c9",x"05",x"ab",x"f0"),
  1679 => (x"c3",x"ec",x"c1",x"87"),
  1680 => (x"c2",x"78",x"c1",x"48"),
  1681 => (x"e0",x"c3",x"87",x"e3"),
  1682 => (x"87",x"c9",x"05",x"ab"),
  1683 => (x"48",x"c7",x"ec",x"c1"),
  1684 => (x"d4",x"c2",x"78",x"c1"),
  1685 => (x"c7",x"ec",x"c1",x"87"),
  1686 => (x"87",x"c6",x"02",x"bf"),
  1687 => (x"4c",x"a3",x"c0",x"c2"),
  1688 => (x"4c",x"73",x"87",x"c2"),
  1689 => (x"bf",x"c3",x"ec",x"c1"),
  1690 => (x"87",x"e0",x"c0",x"02"),
  1691 => (x"b7",x"c4",x"49",x"74"),
  1692 => (x"ed",x"c1",x"91",x"29"),
  1693 => (x"4a",x"74",x"81",x"da"),
  1694 => (x"92",x"c2",x"9a",x"cf"),
  1695 => (x"30",x"72",x"48",x"c1"),
  1696 => (x"ba",x"ff",x"4a",x"70"),
  1697 => (x"98",x"69",x"48",x"72"),
  1698 => (x"87",x"db",x"79",x"70"),
  1699 => (x"b7",x"c4",x"49",x"74"),
  1700 => (x"ed",x"c1",x"91",x"29"),
  1701 => (x"4a",x"74",x"81",x"da"),
  1702 => (x"92",x"c2",x"9a",x"cf"),
  1703 => (x"30",x"72",x"48",x"c3"),
  1704 => (x"69",x"48",x"4a",x"70"),
  1705 => (x"75",x"79",x"70",x"b0"),
  1706 => (x"f0",x"c0",x"05",x"9d"),
  1707 => (x"48",x"d0",x"ff",x"87"),
  1708 => (x"ff",x"78",x"e1",x"c8"),
  1709 => (x"78",x"c5",x"48",x"d4"),
  1710 => (x"bf",x"c7",x"ec",x"c1"),
  1711 => (x"c3",x"87",x"c3",x"02"),
  1712 => (x"ec",x"c1",x"78",x"e0"),
  1713 => (x"c6",x"02",x"bf",x"c3"),
  1714 => (x"48",x"d4",x"ff",x"87"),
  1715 => (x"ff",x"78",x"f0",x"c3"),
  1716 => (x"0b",x"7b",x"0b",x"d4"),
  1717 => (x"c8",x"48",x"d0",x"ff"),
  1718 => (x"e0",x"c0",x"78",x"e1"),
  1719 => (x"c7",x"ec",x"c1",x"78"),
  1720 => (x"c1",x"78",x"c0",x"48"),
  1721 => (x"c0",x"48",x"c3",x"ec"),
  1722 => (x"fe",x"ed",x"c2",x"78"),
  1723 => (x"87",x"f2",x"f9",x"49"),
  1724 => (x"b7",x"c0",x"4b",x"70"),
  1725 => (x"fe",x"fc",x"03",x"ab"),
  1726 => (x"26",x"48",x"c0",x"87"),
  1727 => (x"26",x"4c",x"26",x"4d"),
  1728 => (x"00",x"4f",x"26",x"4b"),
  1729 => (x"00",x"00",x"00",x"00"),
  1730 => (x"1e",x"00",x"00",x"00"),
  1731 => (x"49",x"72",x"4a",x"c0"),
  1732 => (x"ed",x"c1",x"91",x"c4"),
  1733 => (x"79",x"c0",x"81",x"da"),
  1734 => (x"b7",x"d0",x"82",x"c1"),
  1735 => (x"87",x"ee",x"04",x"aa"),
  1736 => (x"5e",x"0e",x"4f",x"26"),
  1737 => (x"0e",x"5d",x"5c",x"5b"),
  1738 => (x"e5",x"f8",x"4d",x"71"),
  1739 => (x"c4",x"4a",x"75",x"87"),
  1740 => (x"c1",x"92",x"2a",x"b7"),
  1741 => (x"75",x"82",x"da",x"ed"),
  1742 => (x"c2",x"9c",x"cf",x"4c"),
  1743 => (x"4b",x"49",x"6a",x"94"),
  1744 => (x"9b",x"c3",x"2b",x"74"),
  1745 => (x"30",x"74",x"48",x"c2"),
  1746 => (x"bc",x"ff",x"4c",x"70"),
  1747 => (x"98",x"71",x"48",x"74"),
  1748 => (x"f5",x"f7",x"7a",x"70"),
  1749 => (x"fe",x"48",x"73",x"87"),
  1750 => (x"00",x"00",x"87",x"e1"),
  1751 => (x"00",x"00",x"00",x"00"),
  1752 => (x"00",x"00",x"00",x"00"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"00",x"00",x"00",x"00"),
  1755 => (x"00",x"00",x"00",x"00"),
  1756 => (x"00",x"00",x"00",x"00"),
  1757 => (x"00",x"00",x"00",x"00"),
  1758 => (x"00",x"00",x"00",x"00"),
  1759 => (x"00",x"00",x"00",x"00"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"ff",x"1e",x"00",x"00"),
  1767 => (x"e1",x"c8",x"48",x"d0"),
  1768 => (x"ff",x"48",x"71",x"78"),
  1769 => (x"26",x"78",x"08",x"d4"),
  1770 => (x"d0",x"ff",x"1e",x"4f"),
  1771 => (x"78",x"e1",x"c8",x"48"),
  1772 => (x"d4",x"ff",x"48",x"71"),
  1773 => (x"66",x"c4",x"78",x"08"),
  1774 => (x"08",x"d4",x"ff",x"48"),
  1775 => (x"1e",x"4f",x"26",x"78"),
  1776 => (x"66",x"c4",x"4a",x"71"),
  1777 => (x"49",x"72",x"1e",x"49"),
  1778 => (x"ff",x"87",x"de",x"ff"),
  1779 => (x"e0",x"c0",x"48",x"d0"),
  1780 => (x"4f",x"26",x"26",x"78"),
  1781 => (x"71",x"1e",x"73",x"1e"),
  1782 => (x"49",x"66",x"c8",x"4b"),
  1783 => (x"c1",x"4a",x"73",x"1e"),
  1784 => (x"ff",x"49",x"a2",x"e0"),
  1785 => (x"c4",x"26",x"87",x"d9"),
  1786 => (x"26",x"4d",x"26",x"87"),
  1787 => (x"26",x"4b",x"26",x"4c"),
  1788 => (x"d4",x"ff",x"1e",x"4f"),
  1789 => (x"7a",x"ff",x"c3",x"4a"),
  1790 => (x"c0",x"48",x"d0",x"ff"),
  1791 => (x"7a",x"de",x"78",x"e1"),
  1792 => (x"bf",x"c8",x"ee",x"c2"),
  1793 => (x"c8",x"48",x"49",x"7a"),
  1794 => (x"71",x"7a",x"70",x"28"),
  1795 => (x"70",x"28",x"d0",x"48"),
  1796 => (x"d8",x"48",x"71",x"7a"),
  1797 => (x"ff",x"7a",x"70",x"28"),
  1798 => (x"e0",x"c0",x"48",x"d0"),
  1799 => (x"1e",x"4f",x"26",x"78"),
  1800 => (x"c8",x"48",x"d0",x"ff"),
  1801 => (x"48",x"71",x"78",x"c9"),
  1802 => (x"78",x"08",x"d4",x"ff"),
  1803 => (x"71",x"1e",x"4f",x"26"),
  1804 => (x"87",x"eb",x"49",x"4a"),
  1805 => (x"c8",x"48",x"d0",x"ff"),
  1806 => (x"1e",x"4f",x"26",x"78"),
  1807 => (x"4b",x"71",x"1e",x"73"),
  1808 => (x"bf",x"d8",x"ee",x"c2"),
  1809 => (x"c2",x"87",x"c3",x"02"),
  1810 => (x"d0",x"ff",x"87",x"eb"),
  1811 => (x"78",x"c9",x"c8",x"48"),
  1812 => (x"e0",x"c0",x"48",x"73"),
  1813 => (x"08",x"d4",x"ff",x"b0"),
  1814 => (x"cc",x"ee",x"c2",x"78"),
  1815 => (x"c8",x"78",x"c0",x"48"),
  1816 => (x"87",x"c5",x"02",x"66"),
  1817 => (x"c2",x"49",x"ff",x"c3"),
  1818 => (x"c2",x"49",x"c0",x"87"),
  1819 => (x"cc",x"59",x"d4",x"ee"),
  1820 => (x"87",x"c6",x"02",x"66"),
  1821 => (x"4a",x"d5",x"d5",x"c5"),
  1822 => (x"ff",x"cf",x"87",x"c4"),
  1823 => (x"ee",x"c2",x"4a",x"ff"),
  1824 => (x"ee",x"c2",x"5a",x"d8"),
  1825 => (x"78",x"c1",x"48",x"d8"),
  1826 => (x"4d",x"26",x"87",x"c4"),
  1827 => (x"4b",x"26",x"4c",x"26"),
  1828 => (x"5e",x"0e",x"4f",x"26"),
  1829 => (x"0e",x"5d",x"5c",x"5b"),
  1830 => (x"ee",x"c2",x"4a",x"71"),
  1831 => (x"72",x"4c",x"bf",x"d4"),
  1832 => (x"87",x"cb",x"02",x"9a"),
  1833 => (x"c1",x"91",x"c8",x"49"),
  1834 => (x"71",x"4b",x"f1",x"f0"),
  1835 => (x"c1",x"87",x"c4",x"83"),
  1836 => (x"c0",x"4b",x"f1",x"f4"),
  1837 => (x"74",x"49",x"13",x"4d"),
  1838 => (x"d0",x"ee",x"c2",x"99"),
  1839 => (x"b8",x"71",x"48",x"bf"),
  1840 => (x"78",x"08",x"d4",x"ff"),
  1841 => (x"85",x"2c",x"b7",x"c1"),
  1842 => (x"04",x"ad",x"b7",x"c8"),
  1843 => (x"ee",x"c2",x"87",x"e7"),
  1844 => (x"c8",x"48",x"bf",x"cc"),
  1845 => (x"d0",x"ee",x"c2",x"80"),
  1846 => (x"87",x"ee",x"fe",x"58"),
  1847 => (x"71",x"1e",x"73",x"1e"),
  1848 => (x"9a",x"4a",x"13",x"4b"),
  1849 => (x"72",x"87",x"cb",x"02"),
  1850 => (x"87",x"e6",x"fe",x"49"),
  1851 => (x"05",x"9a",x"4a",x"13"),
  1852 => (x"d9",x"fe",x"87",x"f5"),
  1853 => (x"ee",x"c2",x"1e",x"87"),
  1854 => (x"c2",x"49",x"bf",x"cc"),
  1855 => (x"c1",x"48",x"cc",x"ee"),
  1856 => (x"c0",x"c4",x"78",x"a1"),
  1857 => (x"db",x"03",x"a9",x"b7"),
  1858 => (x"48",x"d4",x"ff",x"87"),
  1859 => (x"bf",x"d0",x"ee",x"c2"),
  1860 => (x"cc",x"ee",x"c2",x"78"),
  1861 => (x"ee",x"c2",x"49",x"bf"),
  1862 => (x"a1",x"c1",x"48",x"cc"),
  1863 => (x"b7",x"c0",x"c4",x"78"),
  1864 => (x"87",x"e5",x"04",x"a9"),
  1865 => (x"c8",x"48",x"d0",x"ff"),
  1866 => (x"d8",x"ee",x"c2",x"78"),
  1867 => (x"26",x"78",x"c0",x"48"),
  1868 => (x"00",x"00",x"00",x"4f"),
  1869 => (x"00",x"00",x"00",x"00"),
  1870 => (x"00",x"00",x"00",x"00"),
  1871 => (x"00",x"00",x"5f",x"5f"),
  1872 => (x"03",x"03",x"00",x"00"),
  1873 => (x"00",x"03",x"03",x"00"),
  1874 => (x"7f",x"7f",x"14",x"00"),
  1875 => (x"14",x"7f",x"7f",x"14"),
  1876 => (x"2e",x"24",x"00",x"00"),
  1877 => (x"12",x"3a",x"6b",x"6b"),
  1878 => (x"36",x"6a",x"4c",x"00"),
  1879 => (x"32",x"56",x"6c",x"18"),
  1880 => (x"4f",x"7e",x"30",x"00"),
  1881 => (x"68",x"3a",x"77",x"59"),
  1882 => (x"04",x"00",x"00",x"40"),
  1883 => (x"00",x"00",x"03",x"07"),
  1884 => (x"1c",x"00",x"00",x"00"),
  1885 => (x"00",x"41",x"63",x"3e"),
  1886 => (x"41",x"00",x"00",x"00"),
  1887 => (x"00",x"1c",x"3e",x"63"),
  1888 => (x"3e",x"2a",x"08",x"00"),
  1889 => (x"2a",x"3e",x"1c",x"1c"),
  1890 => (x"08",x"08",x"00",x"08"),
  1891 => (x"08",x"08",x"3e",x"3e"),
  1892 => (x"80",x"00",x"00",x"00"),
  1893 => (x"00",x"00",x"60",x"e0"),
  1894 => (x"08",x"08",x"00",x"00"),
  1895 => (x"08",x"08",x"08",x"08"),
  1896 => (x"00",x"00",x"00",x"00"),
  1897 => (x"00",x"00",x"60",x"60"),
  1898 => (x"30",x"60",x"40",x"00"),
  1899 => (x"03",x"06",x"0c",x"18"),
  1900 => (x"7f",x"3e",x"00",x"01"),
  1901 => (x"3e",x"7f",x"4d",x"59"),
  1902 => (x"06",x"04",x"00",x"00"),
  1903 => (x"00",x"00",x"7f",x"7f"),
  1904 => (x"63",x"42",x"00",x"00"),
  1905 => (x"46",x"4f",x"59",x"71"),
  1906 => (x"63",x"22",x"00",x"00"),
  1907 => (x"36",x"7f",x"49",x"49"),
  1908 => (x"16",x"1c",x"18",x"00"),
  1909 => (x"10",x"7f",x"7f",x"13"),
  1910 => (x"67",x"27",x"00",x"00"),
  1911 => (x"39",x"7d",x"45",x"45"),
  1912 => (x"7e",x"3c",x"00",x"00"),
  1913 => (x"30",x"79",x"49",x"4b"),
  1914 => (x"01",x"01",x"00",x"00"),
  1915 => (x"07",x"0f",x"79",x"71"),
  1916 => (x"7f",x"36",x"00",x"00"),
  1917 => (x"36",x"7f",x"49",x"49"),
  1918 => (x"4f",x"06",x"00",x"00"),
  1919 => (x"1e",x"3f",x"69",x"49"),
  1920 => (x"00",x"00",x"00",x"00"),
  1921 => (x"00",x"00",x"66",x"66"),
  1922 => (x"80",x"00",x"00",x"00"),
  1923 => (x"00",x"00",x"66",x"e6"),
  1924 => (x"08",x"08",x"00",x"00"),
  1925 => (x"22",x"22",x"14",x"14"),
  1926 => (x"14",x"14",x"00",x"00"),
  1927 => (x"14",x"14",x"14",x"14"),
  1928 => (x"22",x"22",x"00",x"00"),
  1929 => (x"08",x"08",x"14",x"14"),
  1930 => (x"03",x"02",x"00",x"00"),
  1931 => (x"06",x"0f",x"59",x"51"),
  1932 => (x"41",x"7f",x"3e",x"00"),
  1933 => (x"1e",x"1f",x"55",x"5d"),
  1934 => (x"7f",x"7e",x"00",x"00"),
  1935 => (x"7e",x"7f",x"09",x"09"),
  1936 => (x"7f",x"7f",x"00",x"00"),
  1937 => (x"36",x"7f",x"49",x"49"),
  1938 => (x"3e",x"1c",x"00",x"00"),
  1939 => (x"41",x"41",x"41",x"63"),
  1940 => (x"7f",x"7f",x"00",x"00"),
  1941 => (x"1c",x"3e",x"63",x"41"),
  1942 => (x"7f",x"7f",x"00",x"00"),
  1943 => (x"41",x"41",x"49",x"49"),
  1944 => (x"7f",x"7f",x"00",x"00"),
  1945 => (x"01",x"01",x"09",x"09"),
  1946 => (x"7f",x"3e",x"00",x"00"),
  1947 => (x"7a",x"7b",x"49",x"41"),
  1948 => (x"7f",x"7f",x"00",x"00"),
  1949 => (x"7f",x"7f",x"08",x"08"),
  1950 => (x"41",x"00",x"00",x"00"),
  1951 => (x"00",x"41",x"7f",x"7f"),
  1952 => (x"60",x"20",x"00",x"00"),
  1953 => (x"3f",x"7f",x"40",x"40"),
  1954 => (x"08",x"7f",x"7f",x"00"),
  1955 => (x"41",x"63",x"36",x"1c"),
  1956 => (x"7f",x"7f",x"00",x"00"),
  1957 => (x"40",x"40",x"40",x"40"),
  1958 => (x"06",x"7f",x"7f",x"00"),
  1959 => (x"7f",x"7f",x"06",x"0c"),
  1960 => (x"06",x"7f",x"7f",x"00"),
  1961 => (x"7f",x"7f",x"18",x"0c"),
  1962 => (x"7f",x"3e",x"00",x"00"),
  1963 => (x"3e",x"7f",x"41",x"41"),
  1964 => (x"7f",x"7f",x"00",x"00"),
  1965 => (x"06",x"0f",x"09",x"09"),
  1966 => (x"41",x"7f",x"3e",x"00"),
  1967 => (x"40",x"7e",x"7f",x"61"),
  1968 => (x"7f",x"7f",x"00",x"00"),
  1969 => (x"66",x"7f",x"19",x"09"),
  1970 => (x"6f",x"26",x"00",x"00"),
  1971 => (x"32",x"7b",x"59",x"4d"),
  1972 => (x"01",x"01",x"00",x"00"),
  1973 => (x"01",x"01",x"7f",x"7f"),
  1974 => (x"7f",x"3f",x"00",x"00"),
  1975 => (x"3f",x"7f",x"40",x"40"),
  1976 => (x"3f",x"0f",x"00",x"00"),
  1977 => (x"0f",x"3f",x"70",x"70"),
  1978 => (x"30",x"7f",x"7f",x"00"),
  1979 => (x"7f",x"7f",x"30",x"18"),
  1980 => (x"36",x"63",x"41",x"00"),
  1981 => (x"63",x"36",x"1c",x"1c"),
  1982 => (x"06",x"03",x"01",x"41"),
  1983 => (x"03",x"06",x"7c",x"7c"),
  1984 => (x"59",x"71",x"61",x"01"),
  1985 => (x"41",x"43",x"47",x"4d"),
  1986 => (x"7f",x"00",x"00",x"00"),
  1987 => (x"00",x"41",x"41",x"7f"),
  1988 => (x"06",x"03",x"01",x"00"),
  1989 => (x"60",x"30",x"18",x"0c"),
  1990 => (x"41",x"00",x"00",x"40"),
  1991 => (x"00",x"7f",x"7f",x"41"),
  1992 => (x"06",x"0c",x"08",x"00"),
  1993 => (x"08",x"0c",x"06",x"03"),
  1994 => (x"80",x"80",x"80",x"00"),
  1995 => (x"80",x"80",x"80",x"80"),
  1996 => (x"00",x"00",x"00",x"00"),
  1997 => (x"00",x"04",x"07",x"03"),
  1998 => (x"74",x"20",x"00",x"00"),
  1999 => (x"78",x"7c",x"54",x"54"),
  2000 => (x"7f",x"7f",x"00",x"00"),
  2001 => (x"38",x"7c",x"44",x"44"),
  2002 => (x"7c",x"38",x"00",x"00"),
  2003 => (x"00",x"44",x"44",x"44"),
  2004 => (x"7c",x"38",x"00",x"00"),
  2005 => (x"7f",x"7f",x"44",x"44"),
  2006 => (x"7c",x"38",x"00",x"00"),
  2007 => (x"18",x"5c",x"54",x"54"),
  2008 => (x"7e",x"04",x"00",x"00"),
  2009 => (x"00",x"05",x"05",x"7f"),
  2010 => (x"bc",x"18",x"00",x"00"),
  2011 => (x"7c",x"fc",x"a4",x"a4"),
  2012 => (x"7f",x"7f",x"00",x"00"),
  2013 => (x"78",x"7c",x"04",x"04"),
  2014 => (x"00",x"00",x"00",x"00"),
  2015 => (x"00",x"40",x"7d",x"3d"),
  2016 => (x"80",x"80",x"00",x"00"),
  2017 => (x"00",x"7d",x"fd",x"80"),
  2018 => (x"7f",x"7f",x"00",x"00"),
  2019 => (x"44",x"6c",x"38",x"10"),
  2020 => (x"00",x"00",x"00",x"00"),
  2021 => (x"00",x"40",x"7f",x"3f"),
  2022 => (x"0c",x"7c",x"7c",x"00"),
  2023 => (x"78",x"7c",x"0c",x"18"),
  2024 => (x"7c",x"7c",x"00",x"00"),
  2025 => (x"78",x"7c",x"04",x"04"),
  2026 => (x"7c",x"38",x"00",x"00"),
  2027 => (x"38",x"7c",x"44",x"44"),
  2028 => (x"fc",x"fc",x"00",x"00"),
  2029 => (x"18",x"3c",x"24",x"24"),
  2030 => (x"3c",x"18",x"00",x"00"),
  2031 => (x"fc",x"fc",x"24",x"24"),
  2032 => (x"7c",x"7c",x"00",x"00"),
  2033 => (x"08",x"0c",x"04",x"04"),
  2034 => (x"5c",x"48",x"00",x"00"),
  2035 => (x"20",x"74",x"54",x"54"),
  2036 => (x"3f",x"04",x"00",x"00"),
  2037 => (x"00",x"44",x"44",x"7f"),
  2038 => (x"7c",x"3c",x"00",x"00"),
  2039 => (x"7c",x"7c",x"40",x"40"),
  2040 => (x"3c",x"1c",x"00",x"00"),
  2041 => (x"1c",x"3c",x"60",x"60"),
  2042 => (x"60",x"7c",x"3c",x"00"),
  2043 => (x"3c",x"7c",x"60",x"30"),
  2044 => (x"38",x"6c",x"44",x"00"),
  2045 => (x"44",x"6c",x"38",x"10"),
  2046 => (x"bc",x"1c",x"00",x"00"),
  2047 => (x"1c",x"3c",x"60",x"e0"),
  2048 => (x"64",x"44",x"00",x"00"),
  2049 => (x"44",x"4c",x"5c",x"74"),
  2050 => (x"08",x"08",x"00",x"00"),
  2051 => (x"41",x"41",x"77",x"3e"),
  2052 => (x"00",x"00",x"00",x"00"),
  2053 => (x"00",x"00",x"7f",x"7f"),
  2054 => (x"41",x"41",x"00",x"00"),
  2055 => (x"08",x"08",x"3e",x"77"),
  2056 => (x"01",x"01",x"02",x"00"),
  2057 => (x"01",x"02",x"02",x"03"),
  2058 => (x"7f",x"7f",x"7f",x"00"),
  2059 => (x"7f",x"7f",x"7f",x"7f"),
  2060 => (x"1c",x"08",x"08",x"00"),
  2061 => (x"7f",x"3e",x"3e",x"1c"),
  2062 => (x"3e",x"7f",x"7f",x"7f"),
  2063 => (x"08",x"1c",x"1c",x"3e"),
  2064 => (x"18",x"10",x"00",x"08"),
  2065 => (x"10",x"18",x"7c",x"7c"),
  2066 => (x"30",x"10",x"00",x"00"),
  2067 => (x"10",x"30",x"7c",x"7c"),
  2068 => (x"60",x"30",x"10",x"00"),
  2069 => (x"06",x"1e",x"78",x"60"),
  2070 => (x"3c",x"66",x"42",x"00"),
  2071 => (x"42",x"66",x"3c",x"18"),
  2072 => (x"6a",x"38",x"78",x"00"),
  2073 => (x"38",x"6c",x"c6",x"c2"),
  2074 => (x"00",x"00",x"60",x"00"),
  2075 => (x"60",x"00",x"00",x"60"),
  2076 => (x"5b",x"5e",x"0e",x"00"),
  2077 => (x"1e",x"0e",x"5d",x"5c"),
  2078 => (x"ee",x"c2",x"4c",x"71"),
  2079 => (x"c0",x"4d",x"bf",x"dd"),
  2080 => (x"74",x"1e",x"c0",x"4b"),
  2081 => (x"87",x"c7",x"02",x"ab"),
  2082 => (x"c0",x"48",x"a6",x"c4"),
  2083 => (x"c4",x"87",x"c5",x"78"),
  2084 => (x"78",x"c1",x"48",x"a6"),
  2085 => (x"73",x"1e",x"66",x"c4"),
  2086 => (x"87",x"df",x"ee",x"49"),
  2087 => (x"e0",x"c0",x"86",x"c8"),
  2088 => (x"87",x"ee",x"ef",x"49"),
  2089 => (x"6a",x"4a",x"a5",x"c4"),
  2090 => (x"87",x"f0",x"f0",x"49"),
  2091 => (x"cb",x"87",x"c6",x"f1"),
  2092 => (x"c8",x"83",x"c1",x"85"),
  2093 => (x"ff",x"04",x"ab",x"b7"),
  2094 => (x"26",x"26",x"87",x"c7"),
  2095 => (x"26",x"4c",x"26",x"4d"),
  2096 => (x"1e",x"4f",x"26",x"4b"),
  2097 => (x"ee",x"c2",x"4a",x"71"),
  2098 => (x"ee",x"c2",x"5a",x"e1"),
  2099 => (x"78",x"c7",x"48",x"e1"),
  2100 => (x"87",x"dd",x"fe",x"49"),
  2101 => (x"73",x"1e",x"4f",x"26"),
  2102 => (x"c0",x"4a",x"71",x"1e"),
  2103 => (x"d3",x"03",x"aa",x"b7"),
  2104 => (x"d8",x"d3",x"c2",x"87"),
  2105 => (x"87",x"c4",x"05",x"bf"),
  2106 => (x"87",x"c2",x"4b",x"c1"),
  2107 => (x"d3",x"c2",x"4b",x"c0"),
  2108 => (x"87",x"c4",x"5b",x"dc"),
  2109 => (x"5a",x"dc",x"d3",x"c2"),
  2110 => (x"bf",x"d8",x"d3",x"c2"),
  2111 => (x"c1",x"9a",x"c1",x"4a"),
  2112 => (x"ec",x"49",x"a2",x"c0"),
  2113 => (x"48",x"fc",x"87",x"e8"),
  2114 => (x"bf",x"d8",x"d3",x"c2"),
  2115 => (x"87",x"ef",x"fe",x"78"),
  2116 => (x"c4",x"4a",x"71",x"1e"),
  2117 => (x"49",x"72",x"1e",x"66"),
  2118 => (x"26",x"87",x"f9",x"ea"),
  2119 => (x"ff",x"1e",x"4f",x"26"),
  2120 => (x"ff",x"c3",x"48",x"d4"),
  2121 => (x"48",x"d0",x"ff",x"78"),
  2122 => (x"ff",x"78",x"e1",x"c0"),
  2123 => (x"78",x"c1",x"48",x"d4"),
  2124 => (x"30",x"c4",x"48",x"71"),
  2125 => (x"78",x"08",x"d4",x"ff"),
  2126 => (x"c0",x"48",x"d0",x"ff"),
  2127 => (x"4f",x"26",x"78",x"e0"),
  2128 => (x"5c",x"5b",x"5e",x"0e"),
  2129 => (x"86",x"f4",x"0e",x"5d"),
  2130 => (x"c0",x"48",x"a6",x"c4"),
  2131 => (x"bf",x"ec",x"4b",x"78"),
  2132 => (x"dd",x"ee",x"c2",x"7e"),
  2133 => (x"bf",x"e8",x"4d",x"bf"),
  2134 => (x"d8",x"d3",x"c2",x"4c"),
  2135 => (x"fe",x"e2",x"49",x"bf"),
  2136 => (x"49",x"ee",x"cb",x"87"),
  2137 => (x"cc",x"87",x"f9",x"cd"),
  2138 => (x"49",x"c7",x"58",x"a6"),
  2139 => (x"70",x"87",x"f3",x"e6"),
  2140 => (x"87",x"c8",x"05",x"98"),
  2141 => (x"99",x"c1",x"49",x"6e"),
  2142 => (x"87",x"c3",x"c1",x"02"),
  2143 => (x"bf",x"ec",x"4b",x"c1"),
  2144 => (x"d8",x"d3",x"c2",x"7e"),
  2145 => (x"d6",x"e2",x"49",x"bf"),
  2146 => (x"49",x"66",x"c8",x"87"),
  2147 => (x"70",x"87",x"dd",x"cd"),
  2148 => (x"87",x"d8",x"02",x"98"),
  2149 => (x"bf",x"c0",x"d3",x"c2"),
  2150 => (x"c2",x"b9",x"c1",x"49"),
  2151 => (x"71",x"59",x"c4",x"d3"),
  2152 => (x"cb",x"87",x"fb",x"fd"),
  2153 => (x"f7",x"cc",x"49",x"ee"),
  2154 => (x"58",x"a6",x"cc",x"87"),
  2155 => (x"f1",x"e5",x"49",x"c7"),
  2156 => (x"05",x"98",x"70",x"87"),
  2157 => (x"6e",x"87",x"c5",x"ff"),
  2158 => (x"05",x"99",x"c1",x"49"),
  2159 => (x"73",x"87",x"fd",x"fe"),
  2160 => (x"87",x"d0",x"02",x"9b"),
  2161 => (x"cd",x"fc",x"49",x"ff"),
  2162 => (x"49",x"da",x"c1",x"87"),
  2163 => (x"c4",x"87",x"d3",x"e5"),
  2164 => (x"78",x"c1",x"48",x"a6"),
  2165 => (x"bf",x"d8",x"d3",x"c2"),
  2166 => (x"87",x"d9",x"c1",x"05"),
  2167 => (x"c8",x"48",x"a6",x"c4"),
  2168 => (x"c2",x"78",x"c0",x"c0"),
  2169 => (x"6e",x"7e",x"c4",x"d3"),
  2170 => (x"6e",x"49",x"bf",x"97"),
  2171 => (x"70",x"80",x"c1",x"48"),
  2172 => (x"ed",x"e4",x"71",x"7e"),
  2173 => (x"02",x"98",x"70",x"87"),
  2174 => (x"66",x"c4",x"87",x"c3"),
  2175 => (x"48",x"66",x"c4",x"b4"),
  2176 => (x"c8",x"28",x"b7",x"c1"),
  2177 => (x"98",x"70",x"58",x"a6"),
  2178 => (x"87",x"db",x"ff",x"05"),
  2179 => (x"e4",x"49",x"fd",x"c3"),
  2180 => (x"fa",x"c3",x"87",x"d0"),
  2181 => (x"87",x"ca",x"e4",x"49"),
  2182 => (x"ff",x"c3",x"49",x"74"),
  2183 => (x"c0",x"1e",x"71",x"99"),
  2184 => (x"87",x"ec",x"fb",x"49"),
  2185 => (x"b7",x"c8",x"49",x"74"),
  2186 => (x"c1",x"1e",x"71",x"29"),
  2187 => (x"87",x"e0",x"fb",x"49"),
  2188 => (x"f4",x"c8",x"86",x"c8"),
  2189 => (x"c3",x"49",x"74",x"87"),
  2190 => (x"b7",x"c8",x"99",x"ff"),
  2191 => (x"74",x"b4",x"71",x"2c"),
  2192 => (x"87",x"df",x"02",x"9c"),
  2193 => (x"bf",x"d4",x"d3",x"c2"),
  2194 => (x"87",x"e0",x"ca",x"49"),
  2195 => (x"c0",x"05",x"98",x"70"),
  2196 => (x"4c",x"c0",x"87",x"c4"),
  2197 => (x"e0",x"c2",x"87",x"d3"),
  2198 => (x"87",x"c4",x"ca",x"49"),
  2199 => (x"58",x"d8",x"d3",x"c2"),
  2200 => (x"c2",x"87",x"c6",x"c0"),
  2201 => (x"c0",x"48",x"d4",x"d3"),
  2202 => (x"c2",x"49",x"74",x"78"),
  2203 => (x"ce",x"c0",x"05",x"99"),
  2204 => (x"49",x"eb",x"c3",x"87"),
  2205 => (x"70",x"87",x"eb",x"e2"),
  2206 => (x"02",x"99",x"c2",x"49"),
  2207 => (x"c1",x"87",x"cf",x"c0"),
  2208 => (x"6e",x"7e",x"a5",x"d8"),
  2209 => (x"c5",x"c0",x"02",x"bf"),
  2210 => (x"49",x"fb",x"4b",x"87"),
  2211 => (x"49",x"74",x"0f",x"73"),
  2212 => (x"c0",x"05",x"99",x"c1"),
  2213 => (x"f4",x"c3",x"87",x"ce"),
  2214 => (x"87",x"c6",x"e2",x"49"),
  2215 => (x"99",x"c2",x"49",x"70"),
  2216 => (x"87",x"cf",x"c0",x"02"),
  2217 => (x"7e",x"a5",x"d8",x"c1"),
  2218 => (x"c0",x"02",x"bf",x"6e"),
  2219 => (x"fa",x"4b",x"87",x"c5"),
  2220 => (x"74",x"0f",x"73",x"49"),
  2221 => (x"05",x"99",x"c8",x"49"),
  2222 => (x"c3",x"87",x"ce",x"c0"),
  2223 => (x"e1",x"e1",x"49",x"f5"),
  2224 => (x"c2",x"49",x"70",x"87"),
  2225 => (x"e5",x"c0",x"02",x"99"),
  2226 => (x"e1",x"ee",x"c2",x"87"),
  2227 => (x"ca",x"c0",x"02",x"bf"),
  2228 => (x"88",x"c1",x"48",x"87"),
  2229 => (x"58",x"e5",x"ee",x"c2"),
  2230 => (x"c1",x"87",x"ce",x"c0"),
  2231 => (x"6a",x"4a",x"a5",x"d8"),
  2232 => (x"87",x"c5",x"c0",x"02"),
  2233 => (x"73",x"49",x"ff",x"4b"),
  2234 => (x"48",x"a6",x"c4",x"0f"),
  2235 => (x"49",x"74",x"78",x"c1"),
  2236 => (x"c0",x"05",x"99",x"c4"),
  2237 => (x"f2",x"c3",x"87",x"ce"),
  2238 => (x"87",x"e6",x"e0",x"49"),
  2239 => (x"99",x"c2",x"49",x"70"),
  2240 => (x"87",x"ec",x"c0",x"02"),
  2241 => (x"bf",x"e1",x"ee",x"c2"),
  2242 => (x"b7",x"c7",x"48",x"7e"),
  2243 => (x"cb",x"c0",x"03",x"a8"),
  2244 => (x"c1",x"48",x"6e",x"87"),
  2245 => (x"e5",x"ee",x"c2",x"80"),
  2246 => (x"87",x"cf",x"c0",x"58"),
  2247 => (x"7e",x"a5",x"d8",x"c1"),
  2248 => (x"c0",x"02",x"bf",x"6e"),
  2249 => (x"fe",x"4b",x"87",x"c5"),
  2250 => (x"c4",x"0f",x"73",x"49"),
  2251 => (x"78",x"c1",x"48",x"a6"),
  2252 => (x"ff",x"49",x"fd",x"c3"),
  2253 => (x"70",x"87",x"eb",x"df"),
  2254 => (x"02",x"99",x"c2",x"49"),
  2255 => (x"c2",x"87",x"e5",x"c0"),
  2256 => (x"02",x"bf",x"e1",x"ee"),
  2257 => (x"c2",x"87",x"c9",x"c0"),
  2258 => (x"c0",x"48",x"e1",x"ee"),
  2259 => (x"87",x"cf",x"c0",x"78"),
  2260 => (x"7e",x"a5",x"d8",x"c1"),
  2261 => (x"c0",x"02",x"bf",x"6e"),
  2262 => (x"fd",x"4b",x"87",x"c5"),
  2263 => (x"c4",x"0f",x"73",x"49"),
  2264 => (x"78",x"c1",x"48",x"a6"),
  2265 => (x"ff",x"49",x"fa",x"c3"),
  2266 => (x"70",x"87",x"f7",x"de"),
  2267 => (x"02",x"99",x"c2",x"49"),
  2268 => (x"c2",x"87",x"e9",x"c0"),
  2269 => (x"48",x"bf",x"e1",x"ee"),
  2270 => (x"03",x"a8",x"b7",x"c7"),
  2271 => (x"c2",x"87",x"c9",x"c0"),
  2272 => (x"c7",x"48",x"e1",x"ee"),
  2273 => (x"87",x"cf",x"c0",x"78"),
  2274 => (x"7e",x"a5",x"d8",x"c1"),
  2275 => (x"c0",x"02",x"bf",x"6e"),
  2276 => (x"fc",x"4b",x"87",x"c5"),
  2277 => (x"c4",x"0f",x"73",x"49"),
  2278 => (x"78",x"c1",x"48",x"a6"),
  2279 => (x"ee",x"c2",x"4b",x"c0"),
  2280 => (x"50",x"c0",x"48",x"dc"),
  2281 => (x"c4",x"49",x"ee",x"cb"),
  2282 => (x"a6",x"cc",x"87",x"f6"),
  2283 => (x"dc",x"ee",x"c2",x"58"),
  2284 => (x"c1",x"05",x"bf",x"97"),
  2285 => (x"49",x"74",x"87",x"de"),
  2286 => (x"05",x"99",x"f0",x"c3"),
  2287 => (x"c1",x"87",x"cd",x"c0"),
  2288 => (x"dd",x"ff",x"49",x"da"),
  2289 => (x"98",x"70",x"87",x"dc"),
  2290 => (x"87",x"c8",x"c1",x"02"),
  2291 => (x"bf",x"e8",x"4b",x"c1"),
  2292 => (x"ff",x"c3",x"49",x"4c"),
  2293 => (x"2c",x"b7",x"c8",x"99"),
  2294 => (x"d3",x"c2",x"b4",x"71"),
  2295 => (x"ff",x"49",x"bf",x"d8"),
  2296 => (x"c8",x"87",x"fc",x"d8"),
  2297 => (x"c3",x"c4",x"49",x"66"),
  2298 => (x"02",x"98",x"70",x"87"),
  2299 => (x"c2",x"87",x"c6",x"c0"),
  2300 => (x"c1",x"48",x"dc",x"ee"),
  2301 => (x"dc",x"ee",x"c2",x"50"),
  2302 => (x"c0",x"05",x"bf",x"97"),
  2303 => (x"49",x"74",x"87",x"d6"),
  2304 => (x"05",x"99",x"f0",x"c3"),
  2305 => (x"c1",x"87",x"c5",x"ff"),
  2306 => (x"dc",x"ff",x"49",x"da"),
  2307 => (x"98",x"70",x"87",x"d4"),
  2308 => (x"87",x"f8",x"fe",x"05"),
  2309 => (x"c0",x"02",x"9b",x"73"),
  2310 => (x"a6",x"c8",x"87",x"dc"),
  2311 => (x"e1",x"ee",x"c2",x"48"),
  2312 => (x"66",x"c8",x"78",x"bf"),
  2313 => (x"75",x"91",x"cb",x"49"),
  2314 => (x"bf",x"6e",x"7e",x"a1"),
  2315 => (x"87",x"c6",x"c0",x"02"),
  2316 => (x"49",x"66",x"c8",x"4b"),
  2317 => (x"66",x"c4",x"0f",x"73"),
  2318 => (x"87",x"c8",x"c0",x"02"),
  2319 => (x"bf",x"e1",x"ee",x"c2"),
  2320 => (x"87",x"ed",x"f0",x"49"),
  2321 => (x"bf",x"dc",x"d3",x"c2"),
  2322 => (x"87",x"dd",x"c0",x"02"),
  2323 => (x"87",x"dc",x"c2",x"49"),
  2324 => (x"c0",x"02",x"98",x"70"),
  2325 => (x"ee",x"c2",x"87",x"d3"),
  2326 => (x"f0",x"49",x"bf",x"e1"),
  2327 => (x"49",x"c0",x"87",x"d3"),
  2328 => (x"c2",x"87",x"f3",x"f1"),
  2329 => (x"c0",x"48",x"dc",x"d3"),
  2330 => (x"f1",x"8e",x"f4",x"78"),
  2331 => (x"5e",x"0e",x"87",x"cd"),
  2332 => (x"0e",x"5d",x"5c",x"5b"),
  2333 => (x"c2",x"4c",x"71",x"1e"),
  2334 => (x"49",x"bf",x"dd",x"ee"),
  2335 => (x"4d",x"a1",x"cd",x"c1"),
  2336 => (x"69",x"81",x"d1",x"c1"),
  2337 => (x"02",x"9c",x"74",x"7e"),
  2338 => (x"a5",x"c4",x"87",x"cf"),
  2339 => (x"c2",x"7b",x"74",x"4b"),
  2340 => (x"49",x"bf",x"dd",x"ee"),
  2341 => (x"6e",x"87",x"ec",x"f0"),
  2342 => (x"05",x"9c",x"74",x"7b"),
  2343 => (x"4b",x"c0",x"87",x"c4"),
  2344 => (x"4b",x"c1",x"87",x"c2"),
  2345 => (x"ed",x"f0",x"49",x"73"),
  2346 => (x"02",x"66",x"d4",x"87"),
  2347 => (x"c0",x"49",x"87",x"c8"),
  2348 => (x"4a",x"70",x"87",x"ee"),
  2349 => (x"4a",x"c0",x"87",x"c2"),
  2350 => (x"5a",x"e0",x"d3",x"c2"),
  2351 => (x"87",x"fb",x"ef",x"26"),
  2352 => (x"00",x"00",x"00",x"00"),
  2353 => (x"14",x"11",x"12",x"58"),
  2354 => (x"23",x"1c",x"1b",x"1d"),
  2355 => (x"94",x"91",x"59",x"5a"),
  2356 => (x"f4",x"eb",x"f2",x"f5"),
  2357 => (x"00",x"00",x"00",x"00"),
  2358 => (x"00",x"00",x"00",x"00"),
  2359 => (x"00",x"00",x"00",x"00"),
  2360 => (x"ff",x"4a",x"71",x"1e"),
  2361 => (x"72",x"49",x"bf",x"c8"),
  2362 => (x"4f",x"26",x"48",x"a1"),
  2363 => (x"bf",x"c8",x"ff",x"1e"),
  2364 => (x"c0",x"c0",x"fe",x"89"),
  2365 => (x"a9",x"c0",x"c0",x"c0"),
  2366 => (x"c0",x"87",x"c4",x"01"),
  2367 => (x"c1",x"87",x"c2",x"4a"),
  2368 => (x"26",x"48",x"72",x"4a"),
  2369 => (x"5b",x"5e",x"0e",x"4f"),
  2370 => (x"71",x"0e",x"5d",x"5c"),
  2371 => (x"4c",x"d4",x"ff",x"4b"),
  2372 => (x"c0",x"48",x"66",x"d0"),
  2373 => (x"ff",x"49",x"d6",x"78"),
  2374 => (x"c3",x"87",x"ff",x"d9"),
  2375 => (x"49",x"6c",x"7c",x"ff"),
  2376 => (x"71",x"99",x"ff",x"c3"),
  2377 => (x"f0",x"c3",x"49",x"4d"),
  2378 => (x"a9",x"e0",x"c1",x"99"),
  2379 => (x"c3",x"87",x"cb",x"05"),
  2380 => (x"48",x"6c",x"7c",x"ff"),
  2381 => (x"66",x"d0",x"98",x"c3"),
  2382 => (x"ff",x"c3",x"78",x"08"),
  2383 => (x"49",x"4a",x"6c",x"7c"),
  2384 => (x"ff",x"c3",x"31",x"c8"),
  2385 => (x"71",x"4a",x"6c",x"7c"),
  2386 => (x"c8",x"49",x"72",x"b2"),
  2387 => (x"7c",x"ff",x"c3",x"31"),
  2388 => (x"b2",x"71",x"4a",x"6c"),
  2389 => (x"31",x"c8",x"49",x"72"),
  2390 => (x"6c",x"7c",x"ff",x"c3"),
  2391 => (x"ff",x"b2",x"71",x"4a"),
  2392 => (x"e0",x"c0",x"48",x"d0"),
  2393 => (x"02",x"9b",x"73",x"78"),
  2394 => (x"7b",x"72",x"87",x"c2"),
  2395 => (x"4d",x"26",x"48",x"75"),
  2396 => (x"4b",x"26",x"4c",x"26"),
  2397 => (x"26",x"1e",x"4f",x"26"),
  2398 => (x"5b",x"5e",x"0e",x"4f"),
  2399 => (x"86",x"f8",x"0e",x"5c"),
  2400 => (x"a6",x"c8",x"1e",x"76"),
  2401 => (x"87",x"fd",x"fd",x"49"),
  2402 => (x"4b",x"70",x"86",x"c4"),
  2403 => (x"a8",x"c2",x"48",x"6e"),
  2404 => (x"87",x"f0",x"c2",x"03"),
  2405 => (x"f0",x"c3",x"4a",x"73"),
  2406 => (x"aa",x"d0",x"c1",x"9a"),
  2407 => (x"c1",x"87",x"c7",x"02"),
  2408 => (x"c2",x"05",x"aa",x"e0"),
  2409 => (x"49",x"73",x"87",x"de"),
  2410 => (x"c3",x"02",x"99",x"c8"),
  2411 => (x"87",x"c6",x"ff",x"87"),
  2412 => (x"9c",x"c3",x"4c",x"73"),
  2413 => (x"c1",x"05",x"ac",x"c2"),
  2414 => (x"66",x"c4",x"87",x"c2"),
  2415 => (x"71",x"31",x"c9",x"49"),
  2416 => (x"4a",x"66",x"c4",x"1e"),
  2417 => (x"ee",x"c2",x"92",x"d4"),
  2418 => (x"81",x"72",x"49",x"e5"),
  2419 => (x"87",x"f7",x"cf",x"fe"),
  2420 => (x"d7",x"ff",x"49",x"d8"),
  2421 => (x"c0",x"c8",x"87",x"c4"),
  2422 => (x"ce",x"dd",x"c2",x"1e"),
  2423 => (x"fd",x"eb",x"fd",x"49"),
  2424 => (x"48",x"d0",x"ff",x"87"),
  2425 => (x"c2",x"78",x"e0",x"c0"),
  2426 => (x"cc",x"1e",x"ce",x"dd"),
  2427 => (x"92",x"d4",x"4a",x"66"),
  2428 => (x"49",x"e5",x"ee",x"c2"),
  2429 => (x"cd",x"fe",x"81",x"72"),
  2430 => (x"86",x"cc",x"87",x"ff"),
  2431 => (x"c1",x"05",x"ac",x"c1"),
  2432 => (x"66",x"c4",x"87",x"c2"),
  2433 => (x"71",x"31",x"c9",x"49"),
  2434 => (x"4a",x"66",x"c4",x"1e"),
  2435 => (x"ee",x"c2",x"92",x"d4"),
  2436 => (x"81",x"72",x"49",x"e5"),
  2437 => (x"87",x"ef",x"ce",x"fe"),
  2438 => (x"1e",x"ce",x"dd",x"c2"),
  2439 => (x"d4",x"4a",x"66",x"c8"),
  2440 => (x"e5",x"ee",x"c2",x"92"),
  2441 => (x"fe",x"81",x"72",x"49"),
  2442 => (x"d7",x"87",x"c0",x"cc"),
  2443 => (x"e9",x"d5",x"ff",x"49"),
  2444 => (x"1e",x"c0",x"c8",x"87"),
  2445 => (x"49",x"ce",x"dd",x"c2"),
  2446 => (x"87",x"fb",x"e9",x"fd"),
  2447 => (x"d0",x"ff",x"86",x"cc"),
  2448 => (x"78",x"e0",x"c0",x"48"),
  2449 => (x"e7",x"fc",x"8e",x"f8"),
  2450 => (x"5b",x"5e",x"0e",x"87"),
  2451 => (x"71",x"0e",x"5d",x"5c"),
  2452 => (x"4c",x"d4",x"ff",x"4a"),
  2453 => (x"c3",x"4d",x"66",x"d0"),
  2454 => (x"c5",x"06",x"ad",x"b7"),
  2455 => (x"c1",x"48",x"c0",x"87"),
  2456 => (x"1e",x"72",x"87",x"e1"),
  2457 => (x"93",x"d4",x"4b",x"75"),
  2458 => (x"83",x"e5",x"ee",x"c2"),
  2459 => (x"c6",x"fe",x"49",x"73"),
  2460 => (x"83",x"c8",x"87",x"c7"),
  2461 => (x"d0",x"ff",x"4b",x"6b"),
  2462 => (x"78",x"e1",x"c8",x"48"),
  2463 => (x"48",x"73",x"7c",x"dd"),
  2464 => (x"70",x"98",x"ff",x"c3"),
  2465 => (x"c8",x"49",x"73",x"7c"),
  2466 => (x"48",x"71",x"29",x"b7"),
  2467 => (x"70",x"98",x"ff",x"c3"),
  2468 => (x"d0",x"49",x"73",x"7c"),
  2469 => (x"48",x"71",x"29",x"b7"),
  2470 => (x"70",x"98",x"ff",x"c3"),
  2471 => (x"d8",x"48",x"73",x"7c"),
  2472 => (x"7c",x"70",x"28",x"b7"),
  2473 => (x"7c",x"7c",x"7c",x"c0"),
  2474 => (x"7c",x"7c",x"7c",x"7c"),
  2475 => (x"7c",x"7c",x"7c",x"7c"),
  2476 => (x"48",x"d0",x"ff",x"7c"),
  2477 => (x"75",x"78",x"e0",x"c0"),
  2478 => (x"ff",x"49",x"dc",x"1e"),
  2479 => (x"c8",x"87",x"c0",x"d4"),
  2480 => (x"fa",x"48",x"73",x"86"),
  2481 => (x"73",x"1e",x"87",x"e8"),
  2482 => (x"1e",x"4b",x"c0",x"1e"),
  2483 => (x"bf",x"c7",x"dc",x"c2"),
  2484 => (x"87",x"f5",x"fd",x"49"),
  2485 => (x"dc",x"c2",x"86",x"c4"),
  2486 => (x"fe",x"49",x"bf",x"cb"),
  2487 => (x"70",x"87",x"d0",x"dd"),
  2488 => (x"87",x"c4",x"05",x"98"),
  2489 => (x"4b",x"f4",x"db",x"c2"),
  2490 => (x"87",x"c4",x"48",x"73"),
  2491 => (x"4c",x"26",x"4d",x"26"),
  2492 => (x"4f",x"26",x"4b",x"26"),
  2493 => (x"20",x"4d",x"4f",x"52"),
  2494 => (x"64",x"61",x"6f",x"6c"),
  2495 => (x"20",x"67",x"6e",x"69"),
  2496 => (x"6c",x"69",x"61",x"66"),
  2497 => (x"0f",x"00",x"64",x"65"),
  2498 => (x"1b",x"00",x"00",x"27"),
  2499 => (x"42",x"00",x"00",x"27"),
  2500 => (x"20",x"20",x"43",x"42"),
  2501 => (x"56",x"20",x"20",x"20"),
  2502 => (x"42",x"00",x"44",x"48"),
  2503 => (x"20",x"20",x"43",x"42"),
  2504 => (x"52",x"20",x"20",x"20"),
  2505 => (x"52",x"00",x"4d",x"4f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

